// Check double frees, over allocation
// Check access to unallocated arrays or elements
// Check push overflow, pop underflow
// Next Message 10000280
`define Reset        1  /* Zero all memory sizes                               */
`define Write        2  /* Write an element                                    */
`define Read         3  /* Read an element                                     */
`define Size         4  /* Size of array                                       */
`define Inc          5  /* Increment size of array if possible                 */
`define Dec          6  /* Decrement size of array if possible                 */
`define Index        7  /* Index of element in array                           */
`define Less         8  /* Elements of array less than in                      */
`define Greater      9  /* Elements of array greater than in                   */
`define Up          10  /* Move array up                                       */
`define Down        11  /* Move array down                                     */
`define Long1       12  /* Move long first step                                */
`define Long2       13  /* Move long last  step                                */
`define Push        14  /* Push if possible                                    */
`define Pop         15  /* Pop if possible                                     */
`define Dump        16  /* Dump                                                */
`define Resize      17  /* Resize an array                                     */
`define Alloc       18  /* Allocate a new array before using it                */
`define Free        19  /* Free an array for reuse                             */
`define Add         20  /* Add to an element returning the new value           */
`define AddAfter    21  /* Add to an element returning the previous value      */
`define Subtract    22  /* Subtract to an element returning the new value      */
`define SubAfter    23  /* Subtract to an element returning the previous value */
`define ShiftLeft   24  /* Shift left                                          */
`define ShiftRight  25  /* Shift right                                         */
`define NotLogical  26  /* Not - logical                                       */
`define Not         27  /* Not - bitwise                                       */
`define Or          28  /* Or                                                  */
`define Xor         29  /* Xor                                                 */
`define And         30  /* And                                                 */

module Memory
#(parameter integer ADDRESS_BITS =  8,                                          // Number of bits in an address
  parameter integer INDEX_BITS   =  3,                                          // Bits in in an index
  parameter integer DATA_BITS    = 16)                                          // Width of an element in bits
 (input wire                    clock,                                          // Clock to drive array operations
  input wire[7:0]               action,                                         // Operation to be performed on array
  input wire [ADDRESS_BITS-1:0] array,                                          // The number of the array to work on
  input wire [INDEX_BITS  -1:0] index,                                          // Index within array
  input wire [DATA_BITS   -1:0] in,                                             // Input data
  output reg [DATA_BITS   -1:0] out,                                            // Output data
  output reg [31:0]             error);                                         // Error

  parameter integer ARRAY_LENGTH = 2**INDEX_BITS;                               // Maximum index
  parameter integer ARRAYS       = 2**ADDRESS_BITS;                             // Number of memory elements for both arrays and elements

  reg [DATA_BITS   -1:0] memory     [ARRAYS-1:0][ARRAY_LENGTH-1:0];             // Memory containing arrays in fixed blocks
  reg [DATA_BITS   -1:0] copy                   [ARRAY_LENGTH-1:0];             // Copy of one array
  reg [INDEX_BITS    :0] arraySizes [ARRAYS-1:0];                               // Current size of each array
  reg [ADDRESS_BITS-1:0] freedArrays[ARRAYS-1:0];                               // Currently freed arrays
  reg                    allocations[ARRAYS-1:0];                               // Currently allocated arrays

  integer allocatedArrays;                                                      // Arrays allocated
  integer freedArraysTop;                                                       // Top of the freed arrays stack
  integer result;                                                               // Result of each array operation
  integer size;                                                                 // Size of current array
  integer moveLongStartArray;                                                   // Source array of move long
  integer moveLongStartIndex;                                                   // Source index of move long
  integer i, a, b;                                                              // Index

  task checkWriteable(input integer err);                                       // Check a memory is writable
    begin
       error = 0;
       if (array >= allocatedArrays) begin
         //$display("Array has not been allocated, array %d", array);
         error = err;
       end
       if (!allocations[array]) begin
         //$display("Array has been freed, array %d", array);
         error = err + 1;
       end
    end
  endtask

  task checkReadable(input integer err);                                        // Check a memory locationis readable
    begin
       checkWriteable(err);
       if (index >= arraySizes[array]) begin
         //$display("Access outside array bounds, array %d, size: %d, access: %d", array, arraySizes[array], index);
         error = err + 2;
       end
    end
  endtask

  task dump;                                                                    // Dump some memory
    begin
      //$display("    %2d %2d %2d", arraySizes[0], arraySizes[1], arraySizes[2]);
      for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
        //$display("%2d  %2d %2d %2d", i, memory[0][i], memory[1][i], memory[2][i]);
      end
      //$display("    %2d %2d %2d", allocations[0], allocations[1], allocations[2]);
    end
  endtask

  always @(posedge clock) begin                                                 // Each transition
    case(action)                                                                // Decode request
      `Reset: begin                                                             // Reset
        freedArraysTop = 0;                                                     // Free all arrays
        allocatedArrays = 0;
      end

      `Write: begin                                                             // Write
        checkWriteable(10000010);
        if (!error) begin
          memory[array][index] = in;
          if (index >= arraySizes[array] && index < ARRAY_LENGTH) begin
            arraySizes[array] = index + 1;
          end
          out = in;
        end
      end

      `Read: begin                                                              // Read
        checkReadable(10000020);
        if (!error) begin
          out = memory[array][index];
        end
      end

      `Size: begin                                                              // Size
        checkWriteable(10000030);
        if (!error) begin
          out = arraySizes[array];
        end
      end

      `Dec: begin                                                               // Decrement
        checkWriteable(10000040);
        if (!error) begin
          if (arraySizes[array] > 0) arraySizes[array] = arraySizes[array] - 1;
          else begin
            //$display("Attempt to decrement empty array, array %d", array); error = 10000044;
          end
        end
      end

      `Inc: begin                                                               // Increment
        checkWriteable(10000050);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;
          else begin
            //$display("Attempt to decrement full array, array %d", array);  error = 10000054;
          end
        end
      end

      `Index: begin                                                             // Index
        checkWriteable(10000060);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] == in) result = i + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Less: begin                                                              // Count less
        checkWriteable(10000070);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] < in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Greater: begin                                                           // Count greater
        checkWriteable(10000080);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] > in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Down: begin                                                              // Down
        checkWriteable(10000270);
        if (!error) begin
          size   = arraySizes[array];
          if (size > 0) begin
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i]; // Copy source array
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                       // Move original array up
              if (i > index && i <= size) begin
                memory[array][i-1] = copy[i];
              end
            end
            out = copy[index];                                                  // Return replaced value
            arraySizes[array] = arraySizes[array] - 1;                          // Decrease array size
          end
          else error = 100000274;                                               // Orignal array was emoty so we cannot shift it down
        end
      end

      `Up: begin                                                                // Up
        checkWriteable(10000090);
        if (!error) begin
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i];   // Copy source array
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Move original array up
            if (i > index && i <= size) begin
              memory[array][i] = copy[i-1];
            end
          end
          memory[array][index] = in;                                            // Insert new value
          if (size < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;   // Increase array size
        end
      end

      `Long1: begin                                                             // Move long start
        checkReadable(10000100);
        if (!error) begin
          moveLongStartArray = array;                                           // Record source
          moveLongStartIndex = index;
        end
      end

      `Long2: begin                                                             // Move long finish
        checkWriteable(10000110);
        if (!error) begin
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Copy from source to target
            if (i < in && index + i < ARRAY_LENGTH && moveLongStartIndex+i < ARRAY_LENGTH) begin
              memory[array][index+i] = memory[moveLongStartArray][moveLongStartIndex+i];
              if (index+i >= arraySizes[array]) arraySizes[array] = index+i+1;
            end
          end
        end
      end

      `Push: begin                                                              // Push
        checkWriteable(10000120);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) begin
            memory[array][arraySizes[array]] = in;
            arraySizes[array] = arraySizes[array] + 1;
          end
          else begin
            //$display("Attempt to push to full array, array %d, value %d", array, in);  error = 10000124;
          end
        end
      end

      `Pop: begin                                                               // Pop
        checkWriteable(10000130);
        if (!error) begin
          if (arraySizes[array] > 0) begin
            arraySizes[array] = arraySizes[array] - 1;
            out = memory[array][arraySizes[array]];
          end
          else begin
            //$display("Attempt to pop empty array, array %d", array); error = 10000134;
          end
        end
      end

      `Dump: begin                                                              // Dump
        dump();
      end

      `Resize: begin                                                            // Resize
        checkWriteable(10000140);
        if (!error) begin
          if (in <= ARRAY_LENGTH) arraySizes[array] = in;
          else begin
            //$display("Attempt to make an array too large, array %d, max %d, size %d", array, ARRAY_LENGTH, in); error = 10000144;
          end
        end
      end

      `Alloc: begin                                                             // Allocate an array
        if (freedArraysTop > 0) begin                                           // Reuse a freed array
          freedArraysTop = freedArraysTop - 1;
          result = freedArrays[freedArraysTop];
        end
        else if (allocatedArrays < ARRAYS-1) begin                              // Allocate a new array - assumes enough memory
          result          = allocatedArrays;
          allocatedArrays = allocatedArrays + 1;
        end
        else begin
          //$display("Out of memory, cannot allocate a new array"); error = 10000270;
        end
        allocations[result] = 1;                                                // Allocated
        arraySizes[result] = 0;                                                 // Empty array
        out = result;
      end

      `Free: begin                                                              // Free an array
        checkWriteable(10000150);
        if (!error) begin
          freedArrays[freedArraysTop] = array;                                  // Relies on the user not re freeing a freed array - we should probably hve another array to prevent this
          allocations[array]          = 0;                                      // No longer allocated
          freedArraysTop = freedArraysTop + 1;
        end
      end

      `Add: begin                                                               // Add to an element
        checkReadable(10000160);
        if (!error) begin
          memory[array][index] = memory[array][index] + in;
          out = memory[array][index];
        end
      end

      `AddAfter: begin                                                          // Add to an element after putting the content of the element on out
        checkReadable(10000170);
        if (!error) begin
        out = memory[array][index];
        memory[array][index] = memory[array][index] + in;
        end
      end

      `Subtract: begin                                                          // Subtract from an element
        checkReadable(10000180);
        if (!error) begin
          memory[array][index] = memory[array][index] - in;
          out = memory[array][index];
        end
      end

      `SubAfter: begin                                                          // Subtract from an element after putting the content of the element on out
        checkReadable(10000190);
        if (!error) begin
          out = memory[array][index];
          memory[array][index] = memory[array][index] - in;
        end
      end

      `ShiftLeft: begin                                                         // Shift left
        checkReadable(10000200);
        if (!error) begin
          memory[array][index] = memory[array][index] << in;
          out = memory[array][index];
        end
      end

      `ShiftRight: begin                                                        // Shift right
        checkReadable(10000210);
        if (!error) begin
          memory[array][index] = memory[array][index] >> in;
          out = memory[array][index];
        end
      end

      `NotLogical: begin                                                        // Not logical
        checkReadable(10000220);
        if (!error) begin
          memory[array][index] = !memory[array][index];
          out = memory[array][index];
        end
      end

      `Not: begin                                                               // Not
        checkReadable(10000230);
        if (!error) begin
          memory[array][index] = ~memory[array][index];
          out = memory[array][index];
        end
      end

      `Or: begin                                                                // Or
        checkReadable(10000240);
        if (!error) begin
          memory[array][index] = memory[array][index] | in;
          out = memory[array][index];
        end
      end

      `Xor: begin                                                               // Xor
        checkReadable(10000250);
        if (!error) begin
          memory[array][index] = memory[array][index] ^ in;
          out = memory[array][index];
        end
      end

      `And: begin                                                               // And
        checkReadable(10000260);
        if (!error) begin
          memory[array][index] = memory[array][index] & in;
          out = memory[array][index];
        end
      end
    endcase
  end
endmodule
//-----------------------------------------------------------------------------
// Fpga test
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga                                                                     // Run test programs
 (input  wire clock,                                                            // Driving clock
  input  wire reset,                                                            // Restart program
  output reg  finished,                                                         // Goes high when the program has finished
  output reg  success);                                                         // Goes high on finish if all the tests passed

  reg                heapClock;                                                 // Clock to drive array operations
  reg [7:0]          heapAction;                                                // Operation to be performed on array
  reg [       9-1:0] heapArray;                                         // The number of the array to work on
  reg [       3-1:0] heapIndex;                                         // Index within array
  reg [      12-1:0] heapIn;                                            // Input data
  reg [      12-1:0] heapOut;                                           // Output data
  reg [31        :0] heapError;                                                 // Error on heap operation if not zero

  Memory                                                                        // Memory module
   #(       9,        3,       12)                          // Address bits, index bits, data bits
    heap(                                                                       // Create heap memory
    .clock  (heapClock),
    .action (heapAction),
    .array  (heapArray),
    .index  (heapIndex),
    .in     (heapIn),
    .out    (heapOut),
    .error  (heapError)
  );
  reg [      12-1:0] localMem[    1165-1:0];                       // Local memory
  reg [      12-1:0]   outMem[      67  -1:0];                       // Out channel
  reg [      12-1:0]    inMem[       1   -1:0];                       // In channel

  integer inMemPos;                                                             // Current position in input channel
  integer outMemPos;                                                            // Position in output channel

  integer ip;                                                                   // Instruction pointer
  integer steps;                                                                // Number of steps executed so far
  integer i, j, k;                                                              // A useful counter

  always @(posedge clock) begin                                                 // Each instruction
    if (reset) begin
      ip             = 0;
      steps          = 0;
      inMemPos       = 0;
      outMemPos      = 0;
      finished       = 0;
      success        = 0;

    end
    else begin
      case(ip)

          0 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1;
        end

          1 :
        begin                                                                   // start
          //$display("AAAA %4d %4d start", steps, ip);
              heapAction = `Reset;                                              // Reset heap memory
              ip = 2;
              heapClock = 1;
        end

          2 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3;
        end

          3 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4;
        end

          4 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 5;
              heapClock = 1;
        end

          5 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 6;
        end

          6 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[0] = heapOut;
              ip = 7;
        end

          7 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 8;
        end

          8 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 9;
        end

          9 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[512] = 3;
              ip = 10;
        end

         10 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 11;
        end

         11 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[512];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 12;
              heapClock = 1;
        end

         12 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 13;
        end

         13 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[513] = 0;
              ip = 14;
        end

         14 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 15;
        end

         15 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[513];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 16;
              heapClock = 1;
        end

         16 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 17;
        end

         17 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[514] = 0;
              ip = 18;
        end

         18 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 19;
        end

         19 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[514];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 20;
              heapClock = 1;
        end

         20 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 21;
        end

         21 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[515] = 0;
              ip = 22;
        end

         22 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 23;
        end

         23 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[515];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 24;
              heapClock = 1;
        end

         24 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 25;
        end

         25 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 26;
        end

         26 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1] = 0;
              ip = 27;
        end

         27 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 28;
        end

         28 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[1] >= 66 ? 4458 : 29;
        end

         29 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[2] = localMem[1] + localMem[1];
              ip = 30;
        end

         30 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 31;
        end

         31 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 32;
              heapClock = 1;
        end

         32 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 33;
        end

         33 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[3] = heapOut;
              ip = 34;
        end

         34 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 35;
        end

         35 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 36;
        end

         36 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 37;
        end

         37 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 38;
        end

         38 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 39;
              heapClock = 1;
        end

         39 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 40;
        end

         40 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[516] = heapOut;                                                     // Data retrieved from heap memory
              ip = 41;
              heapClock = 1;
        end

         41 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 42;
        end

         42 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[4] = localMem[516];
              ip = 43;
        end

         43 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[4] != 0 ? 156 : 44;
        end

         44 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 45;
        end

         45 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 46;
              heapClock = 1;
        end

         46 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 47;
        end

         47 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[5] = heapOut;
              ip = 48;
        end

         48 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 49;
        end

         49 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 50;
        end

         50 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[517] = 1;
              ip = 51;
        end

         51 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 52;
        end

         52 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[517];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 53;
              heapClock = 1;
        end

         53 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 54;
        end

         54 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[518] = 0;
              ip = 55;
        end

         55 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 56;
        end

         56 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[518];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 57;
              heapClock = 1;
        end

         57 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 58;
        end

         58 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 59;
        end

         59 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 60;
              heapClock = 1;
        end

         60 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 61;
        end

         61 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[6] = heapOut;
              ip = 62;
        end

         62 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 63;
        end

         63 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 64;
        end

         64 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[519] = localMem[6];
              ip = 65;
        end

         65 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 66;
        end

         66 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[519];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 67;
              heapClock = 1;
        end

         67 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 68;
        end

         68 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 69;
        end

         69 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 70;
              heapClock = 1;
        end

         70 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 71;
        end

         71 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[7] = heapOut;
              ip = 72;
        end

         72 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 73;
        end

         73 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 74;
        end

         74 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[520] = localMem[7];
              ip = 75;
        end

         75 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 76;
        end

         76 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[520];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 77;
              heapClock = 1;
        end

         77 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 78;
        end

         78 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[521] = 0;
              ip = 79;
        end

         79 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 80;
        end

         80 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[521];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 81;
              heapClock = 1;
        end

         81 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 82;
        end

         82 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[522] = localMem[0];
              ip = 83;
        end

         83 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 84;
        end

         84 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[522];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 85;
              heapClock = 1;
        end

         85 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 86;
        end

         86 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 87;
        end

         87 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 88;
              heapClock = 1;
        end

         88 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 89;
        end

         89 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[523] = heapOut;                                                     // Data retrieved from heap memory
              ip = 90;
              heapClock = 1;
        end

         90 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 91;
        end

         91 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[524] = localMem[523] + 1;
              ip = 92;
        end

         92 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 93;
        end

         93 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[524];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 94;
              heapClock = 1;
        end

         94 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 95;
        end

         95 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 96;
        end

         96 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 97;
              heapClock = 1;
        end

         97 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 98;
        end

         98 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[525] = heapOut;                                                     // Data retrieved from heap memory
              ip = 99;
              heapClock = 1;
        end

         99 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 100;
        end

        100 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[526] = localMem[525];
              ip = 101;
        end

        101 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 102;
        end

        102 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[526];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 103;
              heapClock = 1;
        end

        103 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 104;
        end

        104 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 105;
        end

        105 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 106;
              heapClock = 1;
        end

        106 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 107;
        end

        107 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[527] = heapOut;                                                     // Data retrieved from heap memory
              ip = 108;
              heapClock = 1;
        end

        108 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 109;
        end

        109 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[8] = localMem[527];
              ip = 110;
        end

        110 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[528] = localMem[1];
              ip = 111;
        end

        111 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 112;
        end

        112 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[8];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[528];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 113;
              heapClock = 1;
        end

        113 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 114;
        end

        114 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 115;
        end

        115 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 116;
              heapClock = 1;
        end

        116 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 117;
        end

        117 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[529] = heapOut;                                                     // Data retrieved from heap memory
              ip = 118;
              heapClock = 1;
        end

        118 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 119;
        end

        119 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[9] = localMem[529];
              ip = 120;
        end

        120 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[530] = localMem[2];
              ip = 121;
        end

        121 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 122;
        end

        122 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[9];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[530];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 123;
              heapClock = 1;
        end

        123 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 124;
        end

        124 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 125;
        end

        125 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 126;
              heapClock = 1;
        end

        126 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 127;
        end

        127 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[531] = heapOut;                                                     // Data retrieved from heap memory
              ip = 128;
              heapClock = 1;
        end

        128 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 129;
        end

        129 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[532] = localMem[531] + 1;
              ip = 130;
        end

        130 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 131;
        end

        131 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[532];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 132;
              heapClock = 1;
        end

        132 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 133;
        end

        133 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[533] = localMem[5];
              ip = 134;
        end

        134 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 135;
        end

        135 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[533];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 136;
              heapClock = 1;
        end

        136 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 137;
        end

        137 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 138;
        end

        138 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 139;
              heapClock = 1;
        end

        139 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 140;
        end

        140 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[534] = heapOut;                                                     // Data retrieved from heap memory
              ip = 141;
              heapClock = 1;
        end

        141 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 142;
        end

        142 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[10] = localMem[534];
              ip = 143;
        end

        143 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 144;
        end

        144 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[10];
              ip = 145;
              heapClock = 1;
        end

        145 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 146;
        end

        146 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 147;
        end

        147 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 148;
              heapClock = 1;
        end

        148 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 149;
        end

        149 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[535] = heapOut;                                                     // Data retrieved from heap memory
              ip = 150;
              heapClock = 1;
        end

        150 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 151;
        end

        151 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[11] = localMem[535];
              ip = 152;
        end

        152 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 153;
        end

        153 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[11];
              ip = 154;
              heapClock = 1;
        end

        154 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 155;
        end

        155 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4453;
        end

        156 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 157;
        end

        157 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 158;
        end

        158 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 159;
              heapClock = 1;
        end

        159 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 160;
        end

        160 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[536] = heapOut;                                                     // Data retrieved from heap memory
              ip = 161;
              heapClock = 1;
        end

        161 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 162;
        end

        162 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[12] = localMem[536];
              ip = 163;
        end

        163 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 164;
        end

        164 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 165;
              heapClock = 1;
        end

        165 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 166;
        end

        166 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[537] = heapOut;                                                     // Data retrieved from heap memory
              ip = 167;
              heapClock = 1;
        end

        167 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 168;
        end

        168 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[13] = localMem[537];
              ip = 169;
        end

        169 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[12] >= localMem[13] ? 309 : 170;
        end

        170 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 171;
        end

        171 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 172;
              heapClock = 1;
        end

        172 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 173;
        end

        173 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[538] = heapOut;                                                     // Data retrieved from heap memory
              ip = 174;
              heapClock = 1;
        end

        174 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 175;
        end

        175 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[14] = localMem[538];
              ip = 176;
        end

        176 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[14] != 0 ? 308 : 177;
        end

        177 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 178;
        end

        178 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 179;
              heapClock = 1;
        end

        179 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 180;
        end

        180 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[539] = heapOut;                                                     // Data retrieved from heap memory
              ip = 181;
              heapClock = 1;
        end

        181 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 182;
        end

        182 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[15] = !localMem[539];
              ip = 183;
        end

        183 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[15] == 0 ? 307 : 184;
        end

        184 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 185;
        end

        185 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 186;
              heapClock = 1;
        end

        186 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 187;
        end

        187 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[540] = heapOut;                                                     // Data retrieved from heap memory
              ip = 188;
              heapClock = 1;
        end

        188 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 189;
        end

        189 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[16] = localMem[540];
              ip = 190;
        end

        190 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 191;
        end

        191 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[1];
              heapAction = `Index;
              heapArray  = localMem[16];
              ip = 192;
              heapClock = 1;
        end

        192 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 193;
        end

        193 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[17] = heapOut;
              ip = 194;
        end

        194 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 195;
        end

        195 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 196;
        end

        196 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[17] == 0 ? 209 : 197;
        end

        197 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   197");
        end

        198 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   198");
        end

        199 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   199");
        end

        200 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   200");
        end

        201 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   201");
        end

        202 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   202");
        end

        203 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   203");
        end

        204 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   204");
        end

        205 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   205");
        end

        206 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   206");
        end

        207 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   207");
        end

        208 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   208");
        end

        209 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 210;
        end

        210 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 211;
        end

        211 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[12];
              heapArray  = localMem[16];
              ip = 212;
              heapClock = 1;
        end

        212 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 213;
        end

        213 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 214;
        end

        214 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 215;
              heapClock = 1;
        end

        215 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 216;
        end

        216 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[543] = heapOut;                                                     // Data retrieved from heap memory
              ip = 217;
              heapClock = 1;
        end

        217 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 218;
        end

        218 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[19] = localMem[543];
              ip = 219;
        end

        219 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 220;
        end

        220 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[12];
              heapArray  = localMem[19];
              ip = 221;
              heapClock = 1;
        end

        221 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 222;
        end

        222 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 223;
        end

        223 :
        begin                                                                   // arrayCountGreater
          //$display("AAAA %4d %4d arrayCountGreater", steps, ip);
              heapIn     = localMem[1];
              heapAction = `Greater;
              heapArray  = localMem[16];
              ip = 224;
              heapClock = 1;
        end

        224 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 225;
        end

        225 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[20] = heapOut;
              ip = 226;
        end

        226 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 227;
        end

        227 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 228;
        end

        228 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[20] != 0 ? 263 : 229;
        end

        229 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 230;
        end

        230 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 231;
              heapClock = 1;
        end

        231 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 232;
        end

        232 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[544] = heapOut;                                                     // Data retrieved from heap memory
              ip = 233;
              heapClock = 1;
        end

        233 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 234;
        end

        234 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[21] = localMem[544];
              ip = 235;
        end

        235 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[545] = localMem[1];
              ip = 236;
        end

        236 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 237;
        end

        237 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[21];                                                // Array to write to
              heapIndex   = localMem[12];                                                // Index of element to write to
              heapIn      = localMem[545];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 238;
              heapClock = 1;
        end

        238 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 239;
        end

        239 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 240;
        end

        240 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 241;
              heapClock = 1;
        end

        241 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 242;
        end

        242 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[546] = heapOut;                                                     // Data retrieved from heap memory
              ip = 243;
              heapClock = 1;
        end

        243 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 244;
        end

        244 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[22] = localMem[546];
              ip = 245;
        end

        245 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[547] = localMem[2];
              ip = 246;
        end

        246 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 247;
        end

        247 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[22];                                                // Array to write to
              heapIndex   = localMem[12];                                                // Index of element to write to
              heapIn      = localMem[547];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 248;
              heapClock = 1;
        end

        248 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 249;
        end

        249 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[548] = localMem[12] + 1;
              ip = 250;
        end

        250 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 251;
        end

        251 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[4];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[548];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 252;
              heapClock = 1;
        end

        252 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 253;
        end

        253 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 254;
        end

        254 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 255;
              heapClock = 1;
        end

        255 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 256;
        end

        256 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[549] = heapOut;                                                     // Data retrieved from heap memory
              ip = 257;
              heapClock = 1;
        end

        257 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 258;
        end

        258 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[550] = localMem[549] + 1;
              ip = 259;
        end

        259 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 260;
        end

        260 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[550];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 261;
              heapClock = 1;
        end

        261 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 262;
        end

        262 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4453;
        end

        263 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   263");
        end

        264 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   264");
        end

        265 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed   265");
        end

        266 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   266");
        end

        267 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   267");
        end

        268 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   268");
        end

        269 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   269");
        end

        270 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   270");
        end

        271 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   271");
        end

        272 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   272");
        end

        273 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   273");
        end

        274 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   274");
        end

        275 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   275");
        end

        276 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   276");
        end

        277 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   277");
        end

        278 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   278");
        end

        279 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   279");
        end

        280 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   280");
        end

        281 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   281");
        end

        282 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   282");
        end

        283 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   283");
        end

        284 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   284");
        end

        285 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   285");
        end

        286 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   286");
        end

        287 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   287");
        end

        288 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   288");
        end

        289 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   289");
        end

        290 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   290");
        end

        291 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   291");
        end

        292 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   292");
        end

        293 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   293");
        end

        294 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   294");
        end

        295 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   295");
        end

        296 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   296");
        end

        297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   297");
        end

        298 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   298");
        end

        299 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   299");
        end

        300 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   300");
        end

        301 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   301");
        end

        302 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   302");
        end

        303 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   303");
        end

        304 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   304");
        end

        305 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   305");
        end

        306 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   306");
        end

        307 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 308;
        end

        308 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 309;
        end

        309 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 310;
        end

        310 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 311;
        end

        311 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 312;
              heapClock = 1;
        end

        312 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 313;
        end

        313 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[557] = heapOut;                                                     // Data retrieved from heap memory
              ip = 314;
              heapClock = 1;
        end

        314 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 315;
        end

        315 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[26] = localMem[557];
              ip = 316;
        end

        316 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 317;
        end

        317 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 318;
        end

        318 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 319;
              heapClock = 1;
        end

        319 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 320;
        end

        320 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[558] = heapOut;                                                     // Data retrieved from heap memory
              ip = 321;
              heapClock = 1;
        end

        321 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 322;
        end

        322 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[28] = localMem[558];
              ip = 323;
        end

        323 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 324;
        end

        324 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 325;
              heapClock = 1;
        end

        325 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 326;
        end

        326 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[559] = heapOut;                                                     // Data retrieved from heap memory
              ip = 327;
              heapClock = 1;
        end

        327 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 328;
        end

        328 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[29] = localMem[559];
              ip = 329;
        end

        329 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 330;
        end

        330 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 331;
              heapClock = 1;
        end

        331 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 332;
        end

        332 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[560] = heapOut;                                                     // Data retrieved from heap memory
              ip = 333;
              heapClock = 1;
        end

        333 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 334;
        end

        334 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[30] = localMem[560];
              ip = 335;
        end

        335 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[28] <  localMem[30] ? 1287 : 336;
        end

        336 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[31] = localMem[30];
              ip = 337;
        end

        337 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[31] = localMem[31] >> 1;
              ip = 338;
              ip = 338;
        end

        338 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[32] = localMem[31] + 1;
              ip = 339;
        end

        339 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 340;
        end

        340 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 341;
              heapClock = 1;
        end

        341 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 342;
        end

        342 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[561] = heapOut;                                                     // Data retrieved from heap memory
              ip = 343;
              heapClock = 1;
        end

        343 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 344;
        end

        344 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[33] = localMem[561];
              ip = 345;
        end

        345 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[33] == 0 ? 764 : 346;
        end

        346 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   346");
        end

        347 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   347");
        end

        348 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   348");
        end

        349 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   349");
        end

        350 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   350");
        end

        351 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   351");
        end

        352 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   352");
        end

        353 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   353");
        end

        354 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   354");
        end

        355 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   355");
        end

        356 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   356");
        end

        357 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   357");
        end

        358 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   358");
        end

        359 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   359");
        end

        360 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   360");
        end

        361 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   361");
        end

        362 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   362");
        end

        363 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   363");
        end

        364 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   364");
        end

        365 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   365");
        end

        366 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   366");
        end

        367 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   367");
        end

        368 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   368");
        end

        369 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   369");
        end

        370 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   370");
        end

        371 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   371");
        end

        372 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   372");
        end

        373 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   373");
        end

        374 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   374");
        end

        375 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   375");
        end

        376 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   376");
        end

        377 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   377");
        end

        378 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   378");
        end

        379 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   379");
        end

        380 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   380");
        end

        381 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   381");
        end

        382 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   382");
        end

        383 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   383");
        end

        384 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   384");
        end

        385 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   385");
        end

        386 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   386");
        end

        387 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   387");
        end

        388 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   388");
        end

        389 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   389");
        end

        390 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   390");
        end

        391 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   391");
        end

        392 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   392");
        end

        393 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   393");
        end

        394 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   394");
        end

        395 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   395");
        end

        396 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   396");
        end

        397 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   397");
        end

        398 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   398");
        end

        399 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   399");
        end

        400 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   400");
        end

        401 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   401");
        end

        402 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   402");
        end

        403 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   403");
        end

        404 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   404");
        end

        405 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   405");
        end

        406 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   406");
        end

        407 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   407");
        end

        408 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   408");
        end

        409 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   409");
        end

        410 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   410");
        end

        411 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   411");
        end

        412 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   412");
        end

        413 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   413");
        end

        414 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   414");
        end

        415 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   415");
        end

        416 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   416");
        end

        417 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   417");
        end

        418 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   418");
        end

        419 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   419");
        end

        420 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   420");
        end

        421 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   421");
        end

        422 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   422");
        end

        423 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   423");
        end

        424 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   424");
        end

        425 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   425");
        end

        426 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   426");
        end

        427 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   427");
        end

        428 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   428");
        end

        429 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   429");
        end

        430 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   430");
        end

        431 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   431");
        end

        432 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   432");
        end

        433 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   433");
        end

        434 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   434");
        end

        435 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   435");
        end

        436 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   436");
        end

        437 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   437");
        end

        438 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   438");
        end

        439 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   439");
        end

        440 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   440");
        end

        441 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   441");
        end

        442 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   442");
        end

        443 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   443");
        end

        444 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   444");
        end

        445 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   445");
        end

        446 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   446");
        end

        447 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   447");
        end

        448 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   448");
        end

        449 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   449");
        end

        450 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   450");
        end

        451 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   451");
        end

        452 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   452");
        end

        453 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   453");
        end

        454 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   454");
        end

        455 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   455");
        end

        456 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   456");
        end

        457 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   457");
        end

        458 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   458");
        end

        459 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   459");
        end

        460 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   460");
        end

        461 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   461");
        end

        462 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   462");
        end

        463 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   463");
        end

        464 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   464");
        end

        465 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   465");
        end

        466 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   466");
        end

        467 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   467");
        end

        468 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   468");
        end

        469 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   469");
        end

        470 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   470");
        end

        471 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   471");
        end

        472 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   472");
        end

        473 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   473");
        end

        474 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   474");
        end

        475 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   475");
        end

        476 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   476");
        end

        477 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   477");
        end

        478 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   478");
        end

        479 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   479");
        end

        480 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   480");
        end

        481 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   481");
        end

        482 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   482");
        end

        483 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   483");
        end

        484 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   484");
        end

        485 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   485");
        end

        486 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   486");
        end

        487 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   487");
        end

        488 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   488");
        end

        489 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   489");
        end

        490 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   490");
        end

        491 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   491");
        end

        492 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   492");
        end

        493 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   493");
        end

        494 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   494");
        end

        495 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   495");
        end

        496 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   496");
        end

        497 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   497");
        end

        498 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   498");
        end

        499 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   499");
        end

        500 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   500");
        end

        501 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   501");
        end

        502 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   502");
        end

        503 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   503");
        end

        504 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   504");
        end

        505 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   505");
        end

        506 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   506");
        end

        507 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   507");
        end

        508 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   508");
        end

        509 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   509");
        end

        510 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   510");
        end

        511 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   511");
        end

        512 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   512");
        end

        513 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   513");
        end

        514 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   514");
        end

        515 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   515");
        end

        516 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   516");
        end

        517 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   517");
        end

        518 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   518");
        end

        519 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   519");
        end

        520 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   520");
        end

        521 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   521");
        end

        522 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   522");
        end

        523 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   523");
        end

        524 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   524");
        end

        525 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   525");
        end

        526 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   526");
        end

        527 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   527");
        end

        528 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   528");
        end

        529 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   529");
        end

        530 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   530");
        end

        531 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   531");
        end

        532 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   532");
        end

        533 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   533");
        end

        534 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   534");
        end

        535 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   535");
        end

        536 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   536");
        end

        537 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   537");
        end

        538 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   538");
        end

        539 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   539");
        end

        540 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   540");
        end

        541 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   541");
        end

        542 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   542");
        end

        543 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   543");
        end

        544 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   544");
        end

        545 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   545");
        end

        546 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   546");
        end

        547 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   547");
        end

        548 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   548");
        end

        549 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   549");
        end

        550 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   550");
        end

        551 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   551");
        end

        552 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   552");
        end

        553 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   553");
        end

        554 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   554");
        end

        555 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   555");
        end

        556 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   556");
        end

        557 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   557");
        end

        558 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   558");
        end

        559 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   559");
        end

        560 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   560");
        end

        561 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   561");
        end

        562 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   562");
        end

        563 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   563");
        end

        564 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   564");
        end

        565 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   565");
        end

        566 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   566");
        end

        567 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   567");
        end

        568 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   568");
        end

        569 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   569");
        end

        570 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   570");
        end

        571 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   571");
        end

        572 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   572");
        end

        573 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   573");
        end

        574 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   574");
        end

        575 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   575");
        end

        576 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   576");
        end

        577 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   577");
        end

        578 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   578");
        end

        579 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   579");
        end

        580 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   580");
        end

        581 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   581");
        end

        582 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   582");
        end

        583 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   583");
        end

        584 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   584");
        end

        585 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   585");
        end

        586 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   586");
        end

        587 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   587");
        end

        588 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   588");
        end

        589 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   589");
        end

        590 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   590");
        end

        591 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   591");
        end

        592 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   592");
        end

        593 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   593");
        end

        594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   594");
        end

        595 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   595");
        end

        596 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   596");
        end

        597 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   597");
        end

        598 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   598");
        end

        599 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   599");
        end

        600 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   600");
        end

        601 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   601");
        end

        602 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   602");
        end

        603 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   603");
        end

        604 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   604");
        end

        605 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   605");
        end

        606 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   606");
        end

        607 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   607");
        end

        608 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   608");
        end

        609 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   609");
        end

        610 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   610");
        end

        611 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   611");
        end

        612 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   612");
        end

        613 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   613");
        end

        614 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   614");
        end

        615 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   615");
        end

        616 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   616");
        end

        617 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   617");
        end

        618 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   618");
        end

        619 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   619");
        end

        620 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   620");
        end

        621 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   621");
        end

        622 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   622");
        end

        623 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   623");
        end

        624 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   624");
        end

        625 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   625");
        end

        626 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   626");
        end

        627 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   627");
        end

        628 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   628");
        end

        629 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   629");
        end

        630 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   630");
        end

        631 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   631");
        end

        632 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   632");
        end

        633 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   633");
        end

        634 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   634");
        end

        635 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   635");
        end

        636 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   636");
        end

        637 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   637");
        end

        638 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   638");
        end

        639 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   639");
        end

        640 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   640");
        end

        641 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   641");
        end

        642 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   642");
        end

        643 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   643");
        end

        644 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   644");
        end

        645 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   645");
        end

        646 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   646");
        end

        647 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   647");
        end

        648 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   648");
        end

        649 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   649");
        end

        650 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   650");
        end

        651 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   651");
        end

        652 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   652");
        end

        653 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   653");
        end

        654 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   654");
        end

        655 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   655");
        end

        656 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   656");
        end

        657 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   657");
        end

        658 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   658");
        end

        659 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   659");
        end

        660 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   660");
        end

        661 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   661");
        end

        662 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   662");
        end

        663 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   663");
        end

        664 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   664");
        end

        665 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   665");
        end

        666 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   666");
        end

        667 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   667");
        end

        668 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   668");
        end

        669 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   669");
        end

        670 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   670");
        end

        671 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   671");
        end

        672 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   672");
        end

        673 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   673");
        end

        674 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   674");
        end

        675 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   675");
        end

        676 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   676");
        end

        677 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   677");
        end

        678 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   678");
        end

        679 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   679");
        end

        680 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   680");
        end

        681 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   681");
        end

        682 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   682");
        end

        683 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   683");
        end

        684 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   684");
        end

        685 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   685");
        end

        686 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   686");
        end

        687 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   687");
        end

        688 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   688");
        end

        689 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   689");
        end

        690 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   690");
        end

        691 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   691");
        end

        692 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   692");
        end

        693 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   693");
        end

        694 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   694");
        end

        695 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   695");
        end

        696 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   696");
        end

        697 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   697");
        end

        698 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   698");
        end

        699 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   699");
        end

        700 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   700");
        end

        701 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   701");
        end

        702 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   702");
        end

        703 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   703");
        end

        704 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   704");
        end

        705 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   705");
        end

        706 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   706");
        end

        707 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   707");
        end

        708 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   708");
        end

        709 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   709");
        end

        710 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   710");
        end

        711 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   711");
        end

        712 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   712");
        end

        713 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   713");
        end

        714 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   714");
        end

        715 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   715");
        end

        716 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   716");
        end

        717 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   717");
        end

        718 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   718");
        end

        719 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   719");
        end

        720 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   720");
        end

        721 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   721");
        end

        722 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   722");
        end

        723 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   723");
        end

        724 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   724");
        end

        725 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   725");
        end

        726 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   726");
        end

        727 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   727");
        end

        728 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   728");
        end

        729 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   729");
        end

        730 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   730");
        end

        731 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   731");
        end

        732 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   732");
        end

        733 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   733");
        end

        734 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   734");
        end

        735 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   735");
        end

        736 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   736");
        end

        737 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   737");
        end

        738 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   738");
        end

        739 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   739");
        end

        740 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   740");
        end

        741 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   741");
        end

        742 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   742");
        end

        743 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   743");
        end

        744 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   744");
        end

        745 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   745");
        end

        746 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   746");
        end

        747 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   747");
        end

        748 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   748");
        end

        749 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   749");
        end

        750 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   750");
        end

        751 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   751");
        end

        752 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   752");
        end

        753 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   753");
        end

        754 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   754");
        end

        755 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   755");
        end

        756 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   756");
        end

        757 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   757");
        end

        758 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   758");
        end

        759 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   759");
        end

        760 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   760");
        end

        761 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   761");
        end

        762 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   762");
        end

        763 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   763");
        end

        764 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 765;
        end

        765 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 766;
        end

        766 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 767;
              heapClock = 1;
        end

        767 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 768;
        end

        768 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[81] = heapOut;
              ip = 769;
        end

        769 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 770;
        end

        770 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 771;
        end

        771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[619] = localMem[31];
              ip = 772;
        end

        772 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 773;
        end

        773 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[619];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 774;
              heapClock = 1;
        end

        774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 775;
        end

        775 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[620] = 0;
              ip = 776;
        end

        776 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 777;
        end

        777 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[620];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 778;
              heapClock = 1;
        end

        778 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 779;
        end

        779 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 780;
        end

        780 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 781;
              heapClock = 1;
        end

        781 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 782;
        end

        782 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[82] = heapOut;
              ip = 783;
        end

        783 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 784;
        end

        784 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 785;
        end

        785 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[621] = localMem[82];
              ip = 786;
        end

        786 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 787;
        end

        787 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[621];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 788;
              heapClock = 1;
        end

        788 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 789;
        end

        789 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 790;
        end

        790 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 791;
              heapClock = 1;
        end

        791 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 792;
        end

        792 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[83] = heapOut;
              ip = 793;
        end

        793 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 794;
        end

        794 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 795;
        end

        795 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[622] = localMem[83];
              ip = 796;
        end

        796 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 797;
        end

        797 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[622];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 798;
              heapClock = 1;
        end

        798 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 799;
        end

        799 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[623] = 0;
              ip = 800;
        end

        800 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 801;
        end

        801 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[623];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 802;
              heapClock = 1;
        end

        802 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 803;
        end

        803 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[624] = localMem[29];
              ip = 804;
        end

        804 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 805;
        end

        805 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[624];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 806;
              heapClock = 1;
        end

        806 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 807;
        end

        807 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 808;
        end

        808 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 809;
              heapClock = 1;
        end

        809 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 810;
        end

        810 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[625] = heapOut;                                                     // Data retrieved from heap memory
              ip = 811;
              heapClock = 1;
        end

        811 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 812;
        end

        812 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[626] = localMem[625] + 1;
              ip = 813;
        end

        813 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 814;
        end

        814 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[29];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[626];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 815;
              heapClock = 1;
        end

        815 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 816;
        end

        816 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 817;
        end

        817 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 818;
              heapClock = 1;
        end

        818 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 819;
        end

        819 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[627] = heapOut;                                                     // Data retrieved from heap memory
              ip = 820;
              heapClock = 1;
        end

        820 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 821;
        end

        821 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[628] = localMem[627];
              ip = 822;
        end

        822 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 823;
        end

        823 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[628];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 824;
              heapClock = 1;
        end

        824 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 825;
        end

        825 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 826;
        end

        826 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 827;
              heapClock = 1;
        end

        827 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 828;
        end

        828 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[84] = heapOut;
              ip = 829;
        end

        829 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 830;
        end

        830 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 831;
        end

        831 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[629] = localMem[31];
              ip = 832;
        end

        832 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 833;
        end

        833 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[629];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 834;
              heapClock = 1;
        end

        834 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 835;
        end

        835 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[630] = 0;
              ip = 836;
        end

        836 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 837;
        end

        837 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[630];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 838;
              heapClock = 1;
        end

        838 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 839;
        end

        839 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 840;
        end

        840 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 841;
              heapClock = 1;
        end

        841 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 842;
        end

        842 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[85] = heapOut;
              ip = 843;
        end

        843 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 844;
        end

        844 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 845;
        end

        845 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[631] = localMem[85];
              ip = 846;
        end

        846 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 847;
        end

        847 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[631];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 848;
              heapClock = 1;
        end

        848 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 849;
        end

        849 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 850;
        end

        850 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 851;
              heapClock = 1;
        end

        851 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 852;
        end

        852 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[86] = heapOut;
              ip = 853;
        end

        853 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 854;
        end

        854 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 855;
        end

        855 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[632] = localMem[86];
              ip = 856;
        end

        856 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 857;
        end

        857 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[632];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 858;
              heapClock = 1;
        end

        858 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 859;
        end

        859 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[633] = 0;
              ip = 860;
        end

        860 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 861;
        end

        861 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[633];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 862;
              heapClock = 1;
        end

        862 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 863;
        end

        863 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[634] = localMem[29];
              ip = 864;
        end

        864 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 865;
        end

        865 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[634];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 866;
              heapClock = 1;
        end

        866 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 867;
        end

        867 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 868;
        end

        868 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 869;
              heapClock = 1;
        end

        869 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 870;
        end

        870 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[635] = heapOut;                                                     // Data retrieved from heap memory
              ip = 871;
              heapClock = 1;
        end

        871 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 872;
        end

        872 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[636] = localMem[635] + 1;
              ip = 873;
        end

        873 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 874;
        end

        874 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[29];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[636];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 875;
              heapClock = 1;
        end

        875 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 876;
        end

        876 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 877;
        end

        877 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 878;
              heapClock = 1;
        end

        878 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 879;
        end

        879 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[637] = heapOut;                                                     // Data retrieved from heap memory
              ip = 880;
              heapClock = 1;
        end

        880 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 881;
        end

        881 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[638] = localMem[637];
              ip = 882;
        end

        882 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 883;
        end

        883 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[638];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 884;
              heapClock = 1;
        end

        884 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 885;
        end

        885 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 886;
        end

        886 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 887;
              heapClock = 1;
        end

        887 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 888;
        end

        888 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[639] = heapOut;                                                     // Data retrieved from heap memory
              ip = 889;
              heapClock = 1;
        end

        889 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 890;
        end

        890 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[87] = !localMem[639];
              ip = 891;
        end

        891 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[87] != 0 ? 1091 : 892;
        end

        892 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 893;
        end

        893 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 894;
              heapClock = 1;
        end

        894 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 895;
        end

        895 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[88] = heapOut;
              ip = 896;
        end

        896 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 897;
        end

        897 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 898;
        end

        898 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[640] = localMem[88];
              ip = 899;
        end

        899 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 900;
        end

        900 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[640];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 901;
              heapClock = 1;
        end

        901 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 902;
        end

        902 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 903;
        end

        903 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 904;
              heapClock = 1;
        end

        904 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 905;
        end

        905 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[89] = heapOut;
              ip = 906;
        end

        906 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 907;
        end

        907 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 908;
        end

        908 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[641] = localMem[89];
              ip = 909;
        end

        909 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 910;
        end

        910 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[641];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 911;
              heapClock = 1;
        end

        911 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 912;
        end

        912 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 913;
        end

        913 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 914;
              heapClock = 1;
        end

        914 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 915;
        end

        915 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[642] = heapOut;                                                     // Data retrieved from heap memory
              ip = 916;
              heapClock = 1;
        end

        916 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 917;
        end

        917 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[90] = localMem[642];
              ip = 918;
        end

        918 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 919;
        end

        919 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 920;
              heapClock = 1;
        end

        920 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 921;
        end

        921 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[643] = heapOut;                                                     // Data retrieved from heap memory
              ip = 922;
              heapClock = 1;
        end

        922 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 923;
        end

        923 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[91] = localMem[643];
              ip = 924;
        end

        924 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 925;
        end

        925 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 926;
        end

        926 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[90];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 927;
              heapClock = 1;
        end

        927 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 928;
        end

        928 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[91];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 929;
              heapClock = 1;
        end

        929 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 930;
        end

        930 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 931;
        end

        931 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 932;
        end

        932 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 933;
              heapClock = 1;
        end

        933 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 934;
        end

        934 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[644] = heapOut;                                                     // Data retrieved from heap memory
              ip = 935;
              heapClock = 1;
        end

        935 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 936;
        end

        936 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[92] = localMem[644];
              ip = 937;
        end

        937 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 938;
        end

        938 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 939;
              heapClock = 1;
        end

        939 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 940;
        end

        940 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[645] = heapOut;                                                     // Data retrieved from heap memory
              ip = 941;
              heapClock = 1;
        end

        941 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 942;
        end

        942 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[93] = localMem[645];
              ip = 943;
        end

        943 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 944;
        end

        944 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 945;
        end

        945 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[92];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 946;
              heapClock = 1;
        end

        946 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 947;
        end

        947 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[93];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 948;
              heapClock = 1;
        end

        948 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 949;
        end

        949 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 950;
        end

        950 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 951;
        end

        951 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 952;
              heapClock = 1;
        end

        952 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 953;
        end

        953 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[646] = heapOut;                                                     // Data retrieved from heap memory
              ip = 954;
              heapClock = 1;
        end

        954 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 955;
        end

        955 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[94] = localMem[646];
              ip = 956;
        end

        956 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 957;
        end

        957 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 958;
              heapClock = 1;
        end

        958 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 959;
        end

        959 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[647] = heapOut;                                                     // Data retrieved from heap memory
              ip = 960;
              heapClock = 1;
        end

        960 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 961;
        end

        961 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[95] = localMem[647];
              ip = 962;
        end

        962 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[96] = localMem[31] + 1;
              ip = 963;
        end

        963 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 964;
        end

        964 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 965;
        end

        965 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[94];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 966;
              heapClock = 1;
        end

        966 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 967;
        end

        967 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[95];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[96];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 968;
              heapClock = 1;
        end

        968 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 969;
        end

        969 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 970;
        end

        970 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 971;
        end

        971 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 972;
              heapClock = 1;
        end

        972 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 973;
        end

        973 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[648] = heapOut;                                                     // Data retrieved from heap memory
              ip = 974;
              heapClock = 1;
        end

        974 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 975;
        end

        975 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[97] = localMem[648];
              ip = 976;
        end

        976 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 977;
        end

        977 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 978;
              heapClock = 1;
        end

        978 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 979;
        end

        979 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[649] = heapOut;                                                     // Data retrieved from heap memory
              ip = 980;
              heapClock = 1;
        end

        980 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 981;
        end

        981 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[98] = localMem[649];
              ip = 982;
        end

        982 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 983;
        end

        983 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 984;
        end

        984 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[97];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 985;
              heapClock = 1;
        end

        985 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 986;
        end

        986 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[98];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 987;
              heapClock = 1;
        end

        987 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 988;
        end

        988 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 989;
        end

        989 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 990;
        end

        990 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 991;
              heapClock = 1;
        end

        991 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 992;
        end

        992 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[650] = heapOut;                                                     // Data retrieved from heap memory
              ip = 993;
              heapClock = 1;
        end

        993 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 994;
        end

        994 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[99] = localMem[650];
              ip = 995;
        end

        995 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 996;
        end

        996 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 997;
              heapClock = 1;
        end

        997 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 998;
        end

        998 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[651] = heapOut;                                                     // Data retrieved from heap memory
              ip = 999;
              heapClock = 1;
        end

        999 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1000;
        end

       1000 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[100] = localMem[651];
              ip = 1001;
        end

       1001 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1002;
        end

       1002 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1003;
        end

       1003 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[99];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1004;
              heapClock = 1;
        end

       1004 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1005;
        end

       1005 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[100];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1006;
              heapClock = 1;
        end

       1006 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1007;
        end

       1007 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1008;
        end

       1008 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1009;
        end

       1009 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1010;
              heapClock = 1;
        end

       1010 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1011;
        end

       1011 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[652] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1012;
              heapClock = 1;
        end

       1012 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1013;
        end

       1013 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[101] = localMem[652];
              ip = 1014;
        end

       1014 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1015;
        end

       1015 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1016;
              heapClock = 1;
        end

       1016 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1017;
        end

       1017 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[653] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1018;
              heapClock = 1;
        end

       1018 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1019;
        end

       1019 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[102] = localMem[653];
              ip = 1020;
        end

       1020 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[103] = localMem[31] + 1;
              ip = 1021;
        end

       1021 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1022;
        end

       1022 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1023;
        end

       1023 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[101];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1024;
              heapClock = 1;
        end

       1024 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1025;
        end

       1025 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[102];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[103];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1026;
              heapClock = 1;
        end

       1026 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1027;
        end

       1027 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1028;
        end

       1028 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1029;
        end

       1029 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1030;
              heapClock = 1;
        end

       1030 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1031;
        end

       1031 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[654] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1032;
              heapClock = 1;
        end

       1032 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1033;
        end

       1033 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[104] = localMem[654];
              ip = 1034;
        end

       1034 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[105] = localMem[104] + 1;
              ip = 1035;
        end

       1035 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1036;
        end

       1036 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1037;
              heapClock = 1;
        end

       1037 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1038;
        end

       1038 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[655] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1039;
              heapClock = 1;
        end

       1039 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1040;
        end

       1040 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[106] = localMem[655];
              ip = 1041;
        end

       1041 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1042;
        end

       1042 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[107] = 0;
              ip = 1043;
        end

       1043 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1044;
        end

       1044 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[107] >= localMem[105] ? 1058 : 1045;
        end

       1045 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1046;
        end

       1046 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[106];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[107];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1047;
              heapClock = 1;
        end

       1047 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1048;
        end

       1048 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[656] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1049;
              heapClock = 1;
        end

       1049 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1050;
        end

       1050 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[108] = localMem[656];
              ip = 1051;
        end

       1051 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[657] = localMem[81];
              ip = 1052;
        end

       1052 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1053;
        end

       1053 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[108];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[657];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1054;
              heapClock = 1;
        end

       1054 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1055;
        end

       1055 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1056;
        end

       1056 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[107] = localMem[107] + 1;
              ip = 1057;
        end

       1057 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1043;
        end

       1058 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1059;
        end

       1059 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1060;
        end

       1060 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1061;
              heapClock = 1;
        end

       1061 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1062;
        end

       1062 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[658] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1063;
              heapClock = 1;
        end

       1063 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1064;
        end

       1064 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[109] = localMem[658];
              ip = 1065;
        end

       1065 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[110] = localMem[109] + 1;
              ip = 1066;
        end

       1066 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1067;
        end

       1067 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1068;
              heapClock = 1;
        end

       1068 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1069;
        end

       1069 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[659] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1070;
              heapClock = 1;
        end

       1070 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1071;
        end

       1071 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[111] = localMem[659];
              ip = 1072;
        end

       1072 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1073;
        end

       1073 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[112] = 0;
              ip = 1074;
        end

       1074 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1075;
        end

       1075 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[112] >= localMem[110] ? 1089 : 1076;
        end

       1076 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1077;
        end

       1077 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[111];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[112];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1078;
              heapClock = 1;
        end

       1078 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1079;
        end

       1079 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[660] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1080;
              heapClock = 1;
        end

       1080 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1081;
        end

       1081 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[113] = localMem[660];
              ip = 1082;
        end

       1082 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[661] = localMem[84];
              ip = 1083;
        end

       1083 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1084;
        end

       1084 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[113];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[661];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1085;
              heapClock = 1;
        end

       1085 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1086;
        end

       1086 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1087;
        end

       1087 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[112] = localMem[112] + 1;
              ip = 1088;
        end

       1088 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1074;
        end

       1089 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1090;
        end

       1090 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1178;
        end

       1091 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1092;
        end

       1092 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1093;
        end

       1093 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1094;
              heapClock = 1;
        end

       1094 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1095;
        end

       1095 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[114] = heapOut;
              ip = 1096;
        end

       1096 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1097;
        end

       1097 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1098;
        end

       1098 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[662] = localMem[114];
              ip = 1099;
        end

       1099 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1100;
        end

       1100 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[26];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[662];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1101;
              heapClock = 1;
        end

       1101 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1102;
        end

       1102 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1103;
        end

       1103 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1104;
              heapClock = 1;
        end

       1104 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1105;
        end

       1105 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[663] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1106;
              heapClock = 1;
        end

       1106 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1107;
        end

       1107 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[115] = localMem[663];
              ip = 1108;
        end

       1108 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1109;
        end

       1109 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1110;
              heapClock = 1;
        end

       1110 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1111;
        end

       1111 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[664] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1112;
              heapClock = 1;
        end

       1112 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1113;
        end

       1113 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[116] = localMem[664];
              ip = 1114;
        end

       1114 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1115;
        end

       1115 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1116;
        end

       1116 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[115];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1117;
              heapClock = 1;
        end

       1117 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1118;
        end

       1118 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[116];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1119;
              heapClock = 1;
        end

       1119 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1120;
        end

       1120 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1121;
        end

       1121 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1122;
        end

       1122 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1123;
              heapClock = 1;
        end

       1123 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1124;
        end

       1124 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[665] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1125;
              heapClock = 1;
        end

       1125 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1126;
        end

       1126 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[117] = localMem[665];
              ip = 1127;
        end

       1127 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1128;
        end

       1128 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1129;
              heapClock = 1;
        end

       1129 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1130;
        end

       1130 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[666] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1131;
              heapClock = 1;
        end

       1131 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1132;
        end

       1132 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[118] = localMem[666];
              ip = 1133;
        end

       1133 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1134;
        end

       1134 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1135;
        end

       1135 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[117];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1136;
              heapClock = 1;
        end

       1136 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1137;
        end

       1137 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[118];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1138;
              heapClock = 1;
        end

       1138 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1139;
        end

       1139 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1140;
        end

       1140 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1141;
        end

       1141 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1142;
              heapClock = 1;
        end

       1142 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1143;
        end

       1143 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[667] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1144;
              heapClock = 1;
        end

       1144 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1145;
        end

       1145 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[119] = localMem[667];
              ip = 1146;
        end

       1146 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1147;
        end

       1147 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1148;
              heapClock = 1;
        end

       1148 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1149;
        end

       1149 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[668] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1150;
              heapClock = 1;
        end

       1150 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1151;
        end

       1151 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[120] = localMem[668];
              ip = 1152;
        end

       1152 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1153;
        end

       1153 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1154;
        end

       1154 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[119];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1155;
              heapClock = 1;
        end

       1155 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1156;
        end

       1156 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[120];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1157;
              heapClock = 1;
        end

       1157 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1158;
        end

       1158 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1159;
        end

       1159 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1160;
        end

       1160 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1161;
              heapClock = 1;
        end

       1161 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1162;
        end

       1162 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[669] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1163;
              heapClock = 1;
        end

       1163 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1164;
        end

       1164 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[121] = localMem[669];
              ip = 1165;
        end

       1165 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1166;
        end

       1166 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1167;
              heapClock = 1;
        end

       1167 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1168;
        end

       1168 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[670] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1169;
              heapClock = 1;
        end

       1169 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1170;
        end

       1170 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[122] = localMem[670];
              ip = 1171;
        end

       1171 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1172;
        end

       1172 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1173;
        end

       1173 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[121];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1174;
              heapClock = 1;
        end

       1174 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1175;
        end

       1175 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[122];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1176;
              heapClock = 1;
        end

       1176 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1177;
        end

       1177 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1178;
        end

       1178 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1179;
        end

       1179 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[671] = localMem[26];
              ip = 1180;
        end

       1180 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1181;
        end

       1181 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[671];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1182;
              heapClock = 1;
        end

       1182 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1183;
        end

       1183 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[672] = localMem[26];
              ip = 1184;
        end

       1184 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1185;
        end

       1185 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[672];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1186;
              heapClock = 1;
        end

       1186 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1187;
        end

       1187 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1188;
        end

       1188 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1189;
              heapClock = 1;
        end

       1189 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1190;
        end

       1190 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[673] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1191;
              heapClock = 1;
        end

       1191 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1192;
        end

       1192 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[123] = localMem[673];
              ip = 1193;
        end

       1193 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1194;
        end

       1194 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[123];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1195;
              heapClock = 1;
        end

       1195 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1196;
        end

       1196 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[674] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1197;
              heapClock = 1;
        end

       1197 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1198;
        end

       1198 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[124] = localMem[674];
              ip = 1199;
        end

       1199 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1200;
        end

       1200 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1201;
              heapClock = 1;
        end

       1201 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1202;
        end

       1202 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[675] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1203;
              heapClock = 1;
        end

       1203 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1204;
        end

       1204 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[125] = localMem[675];
              ip = 1205;
        end

       1205 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1206;
        end

       1206 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[125];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1207;
              heapClock = 1;
        end

       1207 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1208;
        end

       1208 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[676] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1209;
              heapClock = 1;
        end

       1209 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1210;
        end

       1210 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[126] = localMem[676];
              ip = 1211;
        end

       1211 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1212;
        end

       1212 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1213;
              heapClock = 1;
        end

       1213 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1214;
        end

       1214 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[677] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1215;
              heapClock = 1;
        end

       1215 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1216;
        end

       1216 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[127] = localMem[677];
              ip = 1217;
        end

       1217 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[678] = localMem[124];
              ip = 1218;
        end

       1218 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1219;
        end

       1219 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[127];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[678];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1220;
              heapClock = 1;
        end

       1220 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1221;
        end

       1221 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1222;
        end

       1222 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1223;
              heapClock = 1;
        end

       1223 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1224;
        end

       1224 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[679] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1225;
              heapClock = 1;
        end

       1225 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1226;
        end

       1226 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[128] = localMem[679];
              ip = 1227;
        end

       1227 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[680] = localMem[126];
              ip = 1228;
        end

       1228 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1229;
        end

       1229 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[128];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[680];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1230;
              heapClock = 1;
        end

       1230 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1231;
        end

       1231 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1232;
        end

       1232 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1233;
              heapClock = 1;
        end

       1233 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1234;
        end

       1234 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[681] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1235;
              heapClock = 1;
        end

       1235 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1236;
        end

       1236 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[129] = localMem[681];
              ip = 1237;
        end

       1237 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[682] = localMem[81];
              ip = 1238;
        end

       1238 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1239;
        end

       1239 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[129];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[682];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1240;
              heapClock = 1;
        end

       1240 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1241;
        end

       1241 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1242;
        end

       1242 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1243;
              heapClock = 1;
        end

       1243 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1244;
        end

       1244 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[683] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1245;
              heapClock = 1;
        end

       1245 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1246;
        end

       1246 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[130] = localMem[683];
              ip = 1247;
        end

       1247 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[684] = localMem[84];
              ip = 1248;
        end

       1248 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1249;
        end

       1249 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[130];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[684];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1250;
              heapClock = 1;
        end

       1250 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1251;
        end

       1251 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[685] = 1;
              ip = 1252;
        end

       1252 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1253;
        end

       1253 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[26];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[685];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1254;
              heapClock = 1;
        end

       1254 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1255;
        end

       1255 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1256;
        end

       1256 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1257;
              heapClock = 1;
        end

       1257 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1258;
        end

       1258 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[686] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1259;
              heapClock = 1;
        end

       1259 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1260;
        end

       1260 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[131] = localMem[686];
              ip = 1261;
        end

       1261 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1262;
        end

       1262 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[131];
              ip = 1263;
              heapClock = 1;
        end

       1263 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1264;
        end

       1264 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1265;
        end

       1265 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1266;
              heapClock = 1;
        end

       1266 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1267;
        end

       1267 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[687] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1268;
              heapClock = 1;
        end

       1268 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1269;
        end

       1269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[132] = localMem[687];
              ip = 1270;
        end

       1270 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1271;
        end

       1271 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[132];
              ip = 1272;
              heapClock = 1;
        end

       1272 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1273;
        end

       1273 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1274;
        end

       1274 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1275;
              heapClock = 1;
        end

       1275 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1276;
        end

       1276 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[688] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1277;
              heapClock = 1;
        end

       1277 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1278;
        end

       1278 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[133] = localMem[688];
              ip = 1279;
        end

       1279 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1280;
        end

       1280 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 2;
              heapArray  = localMem[133];
              ip = 1281;
              heapClock = 1;
        end

       1281 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1282;
        end

       1282 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1284;
        end

       1283 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1283");
        end

       1284 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1285;
        end

       1285 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[27] = 1;
              ip = 1286;
        end

       1286 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1289;
        end

       1287 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1288;
        end

       1288 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[27] = 0;
              ip = 1289;
        end

       1289 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1290;
        end

       1290 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1291;
        end

       1291 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1292;
        end

       1292 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[134] = 0;
              ip = 1293;
        end

       1293 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1294;
        end

       1294 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[134] >= 99 ? 3373 : 1295;
        end

       1295 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1296;
        end

       1296 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1297;
              heapClock = 1;
        end

       1297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1298;
        end

       1298 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[689] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1299;
              heapClock = 1;
        end

       1299 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1300;
        end

       1300 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[135] = localMem[689];
              ip = 1301;
        end

       1301 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[136] = localMem[135] - 1;
              ip = 1302;
        end

       1302 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1303;
        end

       1303 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1304;
              heapClock = 1;
        end

       1304 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1305;
        end

       1305 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[690] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1306;
              heapClock = 1;
        end

       1306 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1307;
        end

       1307 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[137] = localMem[690];
              ip = 1308;
        end

       1308 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1309;
        end

       1309 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[137];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[136];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1310;
              heapClock = 1;
        end

       1310 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1311;
        end

       1311 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[691] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1312;
              heapClock = 1;
        end

       1312 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1313;
        end

       1313 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[138] = localMem[691];
              ip = 1314;
        end

       1314 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[1] <= localMem[138] ? 2326 : 1315;
        end

       1315 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1316;
        end

       1316 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1317;
              heapClock = 1;
        end

       1317 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1318;
        end

       1318 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[692] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1319;
              heapClock = 1;
        end

       1319 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1320;
        end

       1320 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[139] = !localMem[692];
              ip = 1321;
        end

       1321 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[139] == 0 ? 1335 : 1322;
        end

       1322 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[693] = localMem[26];
              ip = 1323;
        end

       1323 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1324;
        end

       1324 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[693];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1325;
              heapClock = 1;
        end

       1325 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1326;
        end

       1326 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[694] = 2;
              ip = 1327;
        end

       1327 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1328;
        end

       1328 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[694];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1329;
              heapClock = 1;
        end

       1329 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1330;
        end

       1330 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[695] = localMem[135] - 1;
              ip = 1331;
        end

       1331 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1332;
        end

       1332 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[695];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1333;
              heapClock = 1;
        end

       1333 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1334;
        end

       1334 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3377;
        end

       1335 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1336;
        end

       1336 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1337;
        end

       1337 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1338;
              heapClock = 1;
        end

       1338 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1339;
        end

       1339 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[696] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1340;
              heapClock = 1;
        end

       1340 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1341;
        end

       1341 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[140] = localMem[696];
              ip = 1342;
        end

       1342 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1343;
        end

       1343 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[135];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1344;
              heapClock = 1;
        end

       1344 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1345;
        end

       1345 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[697] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1346;
              heapClock = 1;
        end

       1346 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1347;
        end

       1347 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[141] = localMem[697];
              ip = 1348;
        end

       1348 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1349;
        end

       1349 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1350;
        end

       1350 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1351;
              heapClock = 1;
        end

       1351 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1352;
        end

       1352 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[698] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1353;
              heapClock = 1;
        end

       1353 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1354;
        end

       1354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[143] = localMem[698];
              ip = 1355;
        end

       1355 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1356;
        end

       1356 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1357;
              heapClock = 1;
        end

       1357 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1358;
        end

       1358 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[699] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1359;
              heapClock = 1;
        end

       1359 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1360;
        end

       1360 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[144] = localMem[699];
              ip = 1361;
        end

       1361 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1362;
        end

       1362 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1363;
              heapClock = 1;
        end

       1363 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1364;
        end

       1364 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[700] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1365;
              heapClock = 1;
        end

       1365 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1366;
        end

       1366 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[145] = localMem[700];
              ip = 1367;
        end

       1367 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[143] <  localMem[145] ? 2319 : 1368;
        end

       1368 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[146] = localMem[145];
              ip = 1369;
        end

       1369 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[146] = localMem[146] >> 1;
              ip = 1370;
              ip = 1370;
        end

       1370 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[147] = localMem[146] + 1;
              ip = 1371;
        end

       1371 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1372;
        end

       1372 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1373;
              heapClock = 1;
        end

       1373 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1374;
        end

       1374 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[701] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1375;
              heapClock = 1;
        end

       1375 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1376;
        end

       1376 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[148] = localMem[701];
              ip = 1377;
        end

       1377 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[148] == 0 ? 1796 : 1378;
        end

       1378 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1379;
        end

       1379 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1380;
              heapClock = 1;
        end

       1380 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1381;
        end

       1381 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[149] = heapOut;
              ip = 1382;
        end

       1382 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1383;
        end

       1383 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1384;
        end

       1384 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[702] = localMem[146];
              ip = 1385;
        end

       1385 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1386;
        end

       1386 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[702];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1387;
              heapClock = 1;
        end

       1387 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1388;
        end

       1388 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[703] = 0;
              ip = 1389;
        end

       1389 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1390;
        end

       1390 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[703];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1391;
              heapClock = 1;
        end

       1391 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1392;
        end

       1392 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1393;
        end

       1393 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1394;
              heapClock = 1;
        end

       1394 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1395;
        end

       1395 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[150] = heapOut;
              ip = 1396;
        end

       1396 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1397;
        end

       1397 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1398;
        end

       1398 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[704] = localMem[150];
              ip = 1399;
        end

       1399 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1400;
        end

       1400 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[704];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1401;
              heapClock = 1;
        end

       1401 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1402;
        end

       1402 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1403;
        end

       1403 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1404;
              heapClock = 1;
        end

       1404 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1405;
        end

       1405 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[151] = heapOut;
              ip = 1406;
        end

       1406 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1407;
        end

       1407 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1408;
        end

       1408 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[705] = localMem[151];
              ip = 1409;
        end

       1409 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1410;
        end

       1410 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[705];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1411;
              heapClock = 1;
        end

       1411 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1412;
        end

       1412 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[706] = 0;
              ip = 1413;
        end

       1413 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1414;
        end

       1414 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[706];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1415;
              heapClock = 1;
        end

       1415 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1416;
        end

       1416 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[707] = localMem[144];
              ip = 1417;
        end

       1417 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1418;
        end

       1418 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[707];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1419;
              heapClock = 1;
        end

       1419 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1420;
        end

       1420 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1421;
        end

       1421 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1422;
              heapClock = 1;
        end

       1422 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1423;
        end

       1423 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[708] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1424;
              heapClock = 1;
        end

       1424 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1425;
        end

       1425 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[709] = localMem[708] + 1;
              ip = 1426;
        end

       1426 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1427;
        end

       1427 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[144];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[709];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1428;
              heapClock = 1;
        end

       1428 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1429;
        end

       1429 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1430;
        end

       1430 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1431;
              heapClock = 1;
        end

       1431 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1432;
        end

       1432 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[710] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1433;
              heapClock = 1;
        end

       1433 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1434;
        end

       1434 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[711] = localMem[710];
              ip = 1435;
        end

       1435 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1436;
        end

       1436 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[711];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1437;
              heapClock = 1;
        end

       1437 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1438;
        end

       1438 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1439;
        end

       1439 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1440;
              heapClock = 1;
        end

       1440 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1441;
        end

       1441 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[712] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1442;
              heapClock = 1;
        end

       1442 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1443;
        end

       1443 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[152] = !localMem[712];
              ip = 1444;
        end

       1444 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[152] != 0 ? 1554 : 1445;
        end

       1445 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1446;
        end

       1446 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1447;
              heapClock = 1;
        end

       1447 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1448;
        end

       1448 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[153] = heapOut;
              ip = 1449;
        end

       1449 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1450;
        end

       1450 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1451;
        end

       1451 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[713] = localMem[153];
              ip = 1452;
        end

       1452 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1453;
        end

       1453 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[713];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1454;
              heapClock = 1;
        end

       1454 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1455;
        end

       1455 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1456;
        end

       1456 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1457;
              heapClock = 1;
        end

       1457 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1458;
        end

       1458 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[714] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1459;
              heapClock = 1;
        end

       1459 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1460;
        end

       1460 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[154] = localMem[714];
              ip = 1461;
        end

       1461 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1462;
        end

       1462 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1463;
              heapClock = 1;
        end

       1463 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1464;
        end

       1464 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[715] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1465;
              heapClock = 1;
        end

       1465 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1466;
        end

       1466 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[155] = localMem[715];
              ip = 1467;
        end

       1467 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1468;
        end

       1468 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1469;
        end

       1469 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[154];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1470;
              heapClock = 1;
        end

       1470 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1471;
        end

       1471 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[155];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[146];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1472;
              heapClock = 1;
        end

       1472 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1473;
        end

       1473 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1474;
        end

       1474 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1475;
        end

       1475 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1476;
              heapClock = 1;
        end

       1476 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1477;
        end

       1477 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[716] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1478;
              heapClock = 1;
        end

       1478 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1479;
        end

       1479 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[156] = localMem[716];
              ip = 1480;
        end

       1480 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1481;
        end

       1481 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1482;
              heapClock = 1;
        end

       1482 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1483;
        end

       1483 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[717] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1484;
              heapClock = 1;
        end

       1484 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1485;
        end

       1485 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[157] = localMem[717];
              ip = 1486;
        end

       1486 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1487;
        end

       1487 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1488;
        end

       1488 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[156];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1489;
              heapClock = 1;
        end

       1489 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1490;
        end

       1490 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[157];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[146];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1491;
              heapClock = 1;
        end

       1491 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1492;
        end

       1492 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1493;
        end

       1493 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1494;
        end

       1494 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1495;
              heapClock = 1;
        end

       1495 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1496;
        end

       1496 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[718] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1497;
              heapClock = 1;
        end

       1497 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1498;
        end

       1498 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[158] = localMem[718];
              ip = 1499;
        end

       1499 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1500;
        end

       1500 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1501;
              heapClock = 1;
        end

       1501 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1502;
        end

       1502 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[719] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1503;
              heapClock = 1;
        end

       1503 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1504;
        end

       1504 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[159] = localMem[719];
              ip = 1505;
        end

       1505 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[160] = localMem[146] + 1;
              ip = 1506;
        end

       1506 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1507;
        end

       1507 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1508;
        end

       1508 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[158];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1509;
              heapClock = 1;
        end

       1509 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1510;
        end

       1510 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[159];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[160];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1511;
              heapClock = 1;
        end

       1511 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1512;
        end

       1512 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1513;
        end

       1513 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1514;
        end

       1514 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1515;
              heapClock = 1;
        end

       1515 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1516;
        end

       1516 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[720] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1517;
              heapClock = 1;
        end

       1517 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1518;
        end

       1518 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[161] = localMem[720];
              ip = 1519;
        end

       1519 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[162] = localMem[161] + 1;
              ip = 1520;
        end

       1520 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1521;
        end

       1521 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1522;
              heapClock = 1;
        end

       1522 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1523;
        end

       1523 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[721] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1524;
              heapClock = 1;
        end

       1524 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1525;
        end

       1525 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[163] = localMem[721];
              ip = 1526;
        end

       1526 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1527;
        end

       1527 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[164] = 0;
              ip = 1528;
        end

       1528 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1529;
        end

       1529 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[164] >= localMem[162] ? 1543 : 1530;
        end

       1530 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1531;
        end

       1531 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[163];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[164];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1532;
              heapClock = 1;
        end

       1532 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1533;
        end

       1533 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[722] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1534;
              heapClock = 1;
        end

       1534 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1535;
        end

       1535 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[165] = localMem[722];
              ip = 1536;
        end

       1536 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[723] = localMem[149];
              ip = 1537;
        end

       1537 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1538;
        end

       1538 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[165];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[723];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1539;
              heapClock = 1;
        end

       1539 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1540;
        end

       1540 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1541;
        end

       1541 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[164] = localMem[164] + 1;
              ip = 1542;
        end

       1542 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1528;
        end

       1543 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1544;
        end

       1544 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1545;
        end

       1545 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1546;
              heapClock = 1;
        end

       1546 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1547;
        end

       1547 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[724] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1548;
              heapClock = 1;
        end

       1548 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1549;
        end

       1549 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[166] = localMem[724];
              ip = 1550;
        end

       1550 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1551;
        end

       1551 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[147];
              heapArray  = localMem[166];
              ip = 1552;
              heapClock = 1;
        end

       1552 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1553;
        end

       1553 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1593;
        end

       1554 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1554");
        end

       1555 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1555");
        end

       1556 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1556");
        end

       1557 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1557");
        end

       1558 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1558");
        end

       1559 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1559");
        end

       1560 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1560");
        end

       1561 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1561");
        end

       1562 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1562");
        end

       1563 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1563");
        end

       1564 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1564");
        end

       1565 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1565");
        end

       1566 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1566");
        end

       1567 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1567");
        end

       1568 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1568");
        end

       1569 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1569");
        end

       1570 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1570");
        end

       1571 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1571");
        end

       1572 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1572");
        end

       1573 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1573");
        end

       1574 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1574");
        end

       1575 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1575");
        end

       1576 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1576");
        end

       1577 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1577");
        end

       1578 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1578");
        end

       1579 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1579");
        end

       1580 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1580");
        end

       1581 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1581");
        end

       1582 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1582");
        end

       1583 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1583");
        end

       1584 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1584");
        end

       1585 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1585");
        end

       1586 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1586");
        end

       1587 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1587");
        end

       1588 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1588");
        end

       1589 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1589");
        end

       1590 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1590");
        end

       1591 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1591");
        end

       1592 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1592");
        end

       1593 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1594;
        end

       1594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[729] = localMem[146];
              ip = 1595;
        end

       1595 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1596;
        end

       1596 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[141];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[729];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1597;
              heapClock = 1;
        end

       1597 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1598;
        end

       1598 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[730] = localMem[148];
              ip = 1599;
        end

       1599 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1600;
        end

       1600 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[730];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1601;
              heapClock = 1;
        end

       1601 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1602;
        end

       1602 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1603;
        end

       1603 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1604;
              heapClock = 1;
        end

       1604 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1605;
        end

       1605 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[731] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1606;
              heapClock = 1;
        end

       1606 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1607;
        end

       1607 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[171] = localMem[731];
              ip = 1608;
        end

       1608 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1609;
        end

       1609 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1610;
              heapClock = 1;
        end

       1610 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1611;
        end

       1611 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[732] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1612;
              heapClock = 1;
        end

       1612 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1613;
        end

       1613 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[172] = localMem[732];
              ip = 1614;
        end

       1614 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1615;
        end

       1615 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[172];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[171];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1616;
              heapClock = 1;
        end

       1616 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1617;
        end

       1617 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[733] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1618;
              heapClock = 1;
        end

       1618 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1619;
        end

       1619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[173] = localMem[733];
              ip = 1620;
        end

       1620 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[173] != localMem[141] ? 1700 : 1621;
        end

       1621 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1622;
        end

       1622 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1623;
              heapClock = 1;
        end

       1623 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1624;
        end

       1624 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[734] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1625;
              heapClock = 1;
        end

       1625 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1626;
        end

       1626 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[174] = localMem[734];
              ip = 1627;
        end

       1627 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1628;
        end

       1628 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[174];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[146];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1629;
              heapClock = 1;
        end

       1629 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1630;
        end

       1630 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[735] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1631;
              heapClock = 1;
        end

       1631 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1632;
        end

       1632 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[175] = localMem[735];
              ip = 1633;
        end

       1633 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1634;
        end

       1634 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1635;
              heapClock = 1;
        end

       1635 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1636;
        end

       1636 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[736] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1637;
              heapClock = 1;
        end

       1637 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1638;
        end

       1638 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[176] = localMem[736];
              ip = 1639;
        end

       1639 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[737] = localMem[175];
              ip = 1640;
        end

       1640 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1641;
        end

       1641 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[176];                                                // Array to write to
              heapIndex   = localMem[171];                                                // Index of element to write to
              heapIn      = localMem[737];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1642;
              heapClock = 1;
        end

       1642 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1643;
        end

       1643 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1644;
        end

       1644 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1645;
              heapClock = 1;
        end

       1645 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1646;
        end

       1646 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[738] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1647;
              heapClock = 1;
        end

       1647 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1648;
        end

       1648 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[177] = localMem[738];
              ip = 1649;
        end

       1649 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1650;
        end

       1650 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[177];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[146];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1651;
              heapClock = 1;
        end

       1651 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1652;
        end

       1652 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[739] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1653;
              heapClock = 1;
        end

       1653 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1654;
        end

       1654 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[178] = localMem[739];
              ip = 1655;
        end

       1655 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1656;
        end

       1656 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1657;
              heapClock = 1;
        end

       1657 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1658;
        end

       1658 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[740] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1659;
              heapClock = 1;
        end

       1659 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1660;
        end

       1660 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[179] = localMem[740];
              ip = 1661;
        end

       1661 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[741] = localMem[178];
              ip = 1662;
        end

       1662 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1663;
        end

       1663 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[179];                                                // Array to write to
              heapIndex   = localMem[171];                                                // Index of element to write to
              heapIn      = localMem[741];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1664;
              heapClock = 1;
        end

       1664 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1665;
        end

       1665 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1666;
        end

       1666 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1667;
              heapClock = 1;
        end

       1667 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1668;
        end

       1668 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[742] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1669;
              heapClock = 1;
        end

       1669 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1670;
        end

       1670 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[180] = localMem[742];
              ip = 1671;
        end

       1671 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1672;
        end

       1672 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[146];
              heapArray  = localMem[180];
              ip = 1673;
              heapClock = 1;
        end

       1673 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1674;
        end

       1674 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1675;
        end

       1675 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1676;
              heapClock = 1;
        end

       1676 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1677;
        end

       1677 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[743] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1678;
              heapClock = 1;
        end

       1678 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1679;
        end

       1679 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[181] = localMem[743];
              ip = 1680;
        end

       1680 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1681;
        end

       1681 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[146];
              heapArray  = localMem[181];
              ip = 1682;
              heapClock = 1;
        end

       1682 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1683;
        end

       1683 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[182] = localMem[171] + 1;
              ip = 1684;
        end

       1684 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[744] = localMem[182];
              ip = 1685;
        end

       1685 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1686;
        end

       1686 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[148];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[744];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1687;
              heapClock = 1;
        end

       1687 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1688;
        end

       1688 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1689;
        end

       1689 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 1690;
              heapClock = 1;
        end

       1690 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1691;
        end

       1691 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[745] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1692;
              heapClock = 1;
        end

       1692 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1693;
        end

       1693 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[183] = localMem[745];
              ip = 1694;
        end

       1694 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[746] = localMem[149];
              ip = 1695;
        end

       1695 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1696;
        end

       1696 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[183];                                                // Array to write to
              heapIndex   = localMem[182];                                                // Index of element to write to
              heapIn      = localMem[746];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1697;
              heapClock = 1;
        end

       1697 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1698;
        end

       1698 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2316;
        end

       1699 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1699");
        end

       1700 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1700");
        end

       1701 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  1701");
        end

       1702 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1702");
        end

       1703 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1703");
        end

       1704 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1704");
        end

       1705 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1705");
        end

       1706 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1706");
        end

       1707 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1707");
        end

       1708 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1708");
        end

       1709 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1709");
        end

       1710 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1710");
        end

       1711 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1711");
        end

       1712 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1712");
        end

       1713 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1713");
        end

       1714 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1714");
        end

       1715 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1715");
        end

       1716 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1716");
        end

       1717 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1717");
        end

       1718 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1718");
        end

       1719 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1719");
        end

       1720 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1720");
        end

       1721 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1721");
        end

       1722 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1722");
        end

       1723 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1723");
        end

       1724 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1724");
        end

       1725 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1725");
        end

       1726 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1726");
        end

       1727 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1727");
        end

       1728 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1728");
        end

       1729 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1729");
        end

       1730 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1730");
        end

       1731 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1731");
        end

       1732 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1732");
        end

       1733 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1733");
        end

       1734 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1734");
        end

       1735 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1735");
        end

       1736 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1736");
        end

       1737 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1737");
        end

       1738 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1738");
        end

       1739 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1739");
        end

       1740 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1740");
        end

       1741 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1741");
        end

       1742 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1742");
        end

       1743 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1743");
        end

       1744 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1744");
        end

       1745 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1745");
        end

       1746 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1746");
        end

       1747 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1747");
        end

       1748 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1748");
        end

       1749 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1749");
        end

       1750 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1750");
        end

       1751 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1751");
        end

       1752 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1752");
        end

       1753 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1753");
        end

       1754 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1754");
        end

       1755 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1755");
        end

       1756 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1756");
        end

       1757 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1757");
        end

       1758 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1758");
        end

       1759 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1759");
        end

       1760 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1760");
        end

       1761 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1761");
        end

       1762 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1762");
        end

       1763 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1763");
        end

       1764 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1764");
        end

       1765 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1765");
        end

       1766 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1766");
        end

       1767 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1767");
        end

       1768 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1768");
        end

       1769 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1769");
        end

       1770 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1770");
        end

       1771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1771");
        end

       1772 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1772");
        end

       1773 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1773");
        end

       1774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1774");
        end

       1775 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1775");
        end

       1776 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1776");
        end

       1777 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1777");
        end

       1778 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1778");
        end

       1779 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1779");
        end

       1780 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1780");
        end

       1781 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1781");
        end

       1782 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1782");
        end

       1783 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1783");
        end

       1784 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1784");
        end

       1785 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1785");
        end

       1786 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1786");
        end

       1787 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1787");
        end

       1788 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1788");
        end

       1789 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1789");
        end

       1790 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1790");
        end

       1791 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1791");
        end

       1792 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1792");
        end

       1793 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1793");
        end

       1794 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1794");
        end

       1795 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1795");
        end

       1796 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1796");
        end

       1797 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1797");
        end

       1798 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1798");
        end

       1799 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1799");
        end

       1800 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1800");
        end

       1801 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1801");
        end

       1802 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1802");
        end

       1803 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1803");
        end

       1804 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1804");
        end

       1805 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1805");
        end

       1806 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1806");
        end

       1807 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1807");
        end

       1808 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1808");
        end

       1809 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1809");
        end

       1810 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1810");
        end

       1811 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1811");
        end

       1812 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1812");
        end

       1813 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1813");
        end

       1814 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1814");
        end

       1815 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1815");
        end

       1816 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1816");
        end

       1817 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1817");
        end

       1818 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1818");
        end

       1819 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1819");
        end

       1820 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1820");
        end

       1821 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1821");
        end

       1822 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1822");
        end

       1823 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1823");
        end

       1824 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1824");
        end

       1825 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1825");
        end

       1826 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1826");
        end

       1827 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1827");
        end

       1828 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1828");
        end

       1829 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1829");
        end

       1830 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1830");
        end

       1831 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1831");
        end

       1832 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1832");
        end

       1833 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1833");
        end

       1834 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1834");
        end

       1835 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1835");
        end

       1836 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1836");
        end

       1837 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1837");
        end

       1838 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1838");
        end

       1839 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1839");
        end

       1840 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1840");
        end

       1841 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1841");
        end

       1842 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1842");
        end

       1843 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1843");
        end

       1844 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1844");
        end

       1845 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1845");
        end

       1846 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1846");
        end

       1847 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1847");
        end

       1848 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1848");
        end

       1849 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1849");
        end

       1850 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1850");
        end

       1851 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1851");
        end

       1852 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1852");
        end

       1853 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1853");
        end

       1854 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1854");
        end

       1855 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1855");
        end

       1856 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1856");
        end

       1857 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1857");
        end

       1858 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1858");
        end

       1859 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1859");
        end

       1860 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1860");
        end

       1861 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1861");
        end

       1862 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1862");
        end

       1863 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1863");
        end

       1864 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1864");
        end

       1865 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1865");
        end

       1866 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1866");
        end

       1867 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1867");
        end

       1868 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1868");
        end

       1869 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1869");
        end

       1870 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1870");
        end

       1871 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1871");
        end

       1872 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1872");
        end

       1873 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1873");
        end

       1874 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1874");
        end

       1875 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1875");
        end

       1876 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1876");
        end

       1877 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1877");
        end

       1878 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1878");
        end

       1879 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1879");
        end

       1880 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1880");
        end

       1881 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1881");
        end

       1882 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1882");
        end

       1883 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1883");
        end

       1884 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1884");
        end

       1885 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1885");
        end

       1886 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1886");
        end

       1887 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1887");
        end

       1888 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1888");
        end

       1889 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1889");
        end

       1890 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1890");
        end

       1891 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1891");
        end

       1892 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1892");
        end

       1893 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1893");
        end

       1894 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1894");
        end

       1895 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1895");
        end

       1896 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1896");
        end

       1897 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1897");
        end

       1898 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1898");
        end

       1899 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1899");
        end

       1900 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1900");
        end

       1901 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1901");
        end

       1902 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1902");
        end

       1903 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1903");
        end

       1904 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1904");
        end

       1905 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1905");
        end

       1906 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1906");
        end

       1907 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1907");
        end

       1908 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1908");
        end

       1909 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1909");
        end

       1910 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1910");
        end

       1911 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1911");
        end

       1912 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1912");
        end

       1913 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1913");
        end

       1914 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1914");
        end

       1915 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1915");
        end

       1916 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1916");
        end

       1917 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1917");
        end

       1918 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1918");
        end

       1919 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1919");
        end

       1920 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1920");
        end

       1921 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1921");
        end

       1922 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1922");
        end

       1923 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1923");
        end

       1924 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1924");
        end

       1925 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1925");
        end

       1926 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1926");
        end

       1927 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1927");
        end

       1928 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1928");
        end

       1929 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1929");
        end

       1930 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1930");
        end

       1931 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1931");
        end

       1932 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1932");
        end

       1933 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1933");
        end

       1934 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1934");
        end

       1935 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1935");
        end

       1936 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1936");
        end

       1937 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1937");
        end

       1938 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1938");
        end

       1939 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1939");
        end

       1940 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1940");
        end

       1941 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1941");
        end

       1942 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1942");
        end

       1943 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1943");
        end

       1944 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1944");
        end

       1945 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1945");
        end

       1946 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1946");
        end

       1947 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1947");
        end

       1948 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1948");
        end

       1949 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1949");
        end

       1950 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1950");
        end

       1951 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1951");
        end

       1952 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1952");
        end

       1953 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1953");
        end

       1954 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1954");
        end

       1955 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1955");
        end

       1956 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1956");
        end

       1957 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1957");
        end

       1958 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1958");
        end

       1959 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1959");
        end

       1960 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1960");
        end

       1961 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1961");
        end

       1962 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1962");
        end

       1963 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1963");
        end

       1964 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1964");
        end

       1965 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1965");
        end

       1966 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1966");
        end

       1967 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1967");
        end

       1968 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1968");
        end

       1969 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1969");
        end

       1970 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1970");
        end

       1971 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1971");
        end

       1972 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1972");
        end

       1973 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1973");
        end

       1974 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1974");
        end

       1975 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1975");
        end

       1976 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1976");
        end

       1977 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1977");
        end

       1978 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1978");
        end

       1979 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1979");
        end

       1980 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1980");
        end

       1981 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1981");
        end

       1982 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1982");
        end

       1983 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1983");
        end

       1984 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1984");
        end

       1985 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1985");
        end

       1986 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1986");
        end

       1987 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1987");
        end

       1988 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1988");
        end

       1989 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1989");
        end

       1990 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1990");
        end

       1991 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1991");
        end

       1992 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1992");
        end

       1993 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1993");
        end

       1994 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1994");
        end

       1995 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1995");
        end

       1996 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1996");
        end

       1997 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1997");
        end

       1998 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1998");
        end

       1999 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1999");
        end

       2000 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2000");
        end

       2001 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2001");
        end

       2002 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2002");
        end

       2003 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2003");
        end

       2004 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2004");
        end

       2005 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2005");
        end

       2006 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2006");
        end

       2007 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2007");
        end

       2008 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2008");
        end

       2009 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2009");
        end

       2010 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2010");
        end

       2011 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2011");
        end

       2012 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2012");
        end

       2013 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2013");
        end

       2014 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2014");
        end

       2015 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2015");
        end

       2016 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2016");
        end

       2017 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2017");
        end

       2018 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2018");
        end

       2019 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2019");
        end

       2020 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2020");
        end

       2021 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2021");
        end

       2022 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2022");
        end

       2023 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2023");
        end

       2024 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2024");
        end

       2025 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2025");
        end

       2026 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2026");
        end

       2027 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2027");
        end

       2028 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2028");
        end

       2029 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2029");
        end

       2030 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2030");
        end

       2031 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2031");
        end

       2032 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2032");
        end

       2033 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2033");
        end

       2034 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2034");
        end

       2035 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2035");
        end

       2036 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2036");
        end

       2037 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2037");
        end

       2038 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2038");
        end

       2039 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2039");
        end

       2040 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2040");
        end

       2041 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2041");
        end

       2042 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2042");
        end

       2043 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2043");
        end

       2044 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2044");
        end

       2045 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2045");
        end

       2046 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2046");
        end

       2047 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2047");
        end

       2048 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2048");
        end

       2049 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2049");
        end

       2050 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2050");
        end

       2051 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2051");
        end

       2052 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2052");
        end

       2053 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2053");
        end

       2054 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2054");
        end

       2055 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2055");
        end

       2056 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2056");
        end

       2057 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2057");
        end

       2058 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2058");
        end

       2059 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2059");
        end

       2060 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2060");
        end

       2061 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2061");
        end

       2062 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2062");
        end

       2063 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2063");
        end

       2064 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2064");
        end

       2065 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2065");
        end

       2066 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2066");
        end

       2067 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2067");
        end

       2068 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2068");
        end

       2069 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2069");
        end

       2070 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2070");
        end

       2071 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2071");
        end

       2072 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2072");
        end

       2073 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2073");
        end

       2074 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2074");
        end

       2075 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2075");
        end

       2076 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2076");
        end

       2077 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2077");
        end

       2078 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2078");
        end

       2079 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2079");
        end

       2080 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2080");
        end

       2081 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2081");
        end

       2082 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2082");
        end

       2083 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2083");
        end

       2084 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2084");
        end

       2085 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2085");
        end

       2086 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2086");
        end

       2087 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2087");
        end

       2088 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2088");
        end

       2089 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2089");
        end

       2090 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2090");
        end

       2091 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2091");
        end

       2092 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2092");
        end

       2093 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2093");
        end

       2094 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2094");
        end

       2095 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2095");
        end

       2096 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2096");
        end

       2097 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2097");
        end

       2098 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2098");
        end

       2099 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2099");
        end

       2100 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2100");
        end

       2101 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2101");
        end

       2102 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2102");
        end

       2103 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2103");
        end

       2104 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2104");
        end

       2105 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2105");
        end

       2106 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2106");
        end

       2107 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2107");
        end

       2108 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2108");
        end

       2109 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2109");
        end

       2110 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2110");
        end

       2111 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2111");
        end

       2112 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2112");
        end

       2113 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2113");
        end

       2114 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2114");
        end

       2115 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2115");
        end

       2116 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2116");
        end

       2117 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2117");
        end

       2118 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2118");
        end

       2119 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2119");
        end

       2120 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2120");
        end

       2121 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2121");
        end

       2122 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2122");
        end

       2123 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2123");
        end

       2124 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2124");
        end

       2125 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2125");
        end

       2126 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2126");
        end

       2127 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2127");
        end

       2128 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2128");
        end

       2129 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2129");
        end

       2130 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2130");
        end

       2131 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2131");
        end

       2132 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2132");
        end

       2133 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2133");
        end

       2134 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2134");
        end

       2135 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2135");
        end

       2136 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2136");
        end

       2137 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2137");
        end

       2138 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2138");
        end

       2139 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2139");
        end

       2140 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2140");
        end

       2141 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2141");
        end

       2142 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2142");
        end

       2143 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2143");
        end

       2144 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2144");
        end

       2145 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2145");
        end

       2146 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2146");
        end

       2147 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2147");
        end

       2148 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2148");
        end

       2149 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2149");
        end

       2150 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2150");
        end

       2151 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2151");
        end

       2152 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2152");
        end

       2153 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2153");
        end

       2154 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2154");
        end

       2155 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2155");
        end

       2156 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2156");
        end

       2157 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2157");
        end

       2158 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2158");
        end

       2159 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2159");
        end

       2160 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2160");
        end

       2161 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2161");
        end

       2162 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2162");
        end

       2163 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2163");
        end

       2164 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2164");
        end

       2165 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2165");
        end

       2166 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2166");
        end

       2167 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2167");
        end

       2168 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2168");
        end

       2169 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2169");
        end

       2170 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2170");
        end

       2171 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2171");
        end

       2172 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2172");
        end

       2173 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2173");
        end

       2174 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2174");
        end

       2175 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2175");
        end

       2176 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2176");
        end

       2177 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2177");
        end

       2178 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2178");
        end

       2179 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2179");
        end

       2180 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2180");
        end

       2181 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2181");
        end

       2182 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2182");
        end

       2183 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2183");
        end

       2184 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2184");
        end

       2185 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2185");
        end

       2186 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2186");
        end

       2187 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2187");
        end

       2188 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2188");
        end

       2189 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2189");
        end

       2190 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2190");
        end

       2191 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2191");
        end

       2192 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2192");
        end

       2193 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2193");
        end

       2194 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2194");
        end

       2195 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2195");
        end

       2196 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2196");
        end

       2197 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2197");
        end

       2198 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2198");
        end

       2199 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2199");
        end

       2200 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2200");
        end

       2201 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2201");
        end

       2202 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2202");
        end

       2203 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2203");
        end

       2204 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2204");
        end

       2205 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2205");
        end

       2206 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2206");
        end

       2207 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2207");
        end

       2208 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2208");
        end

       2209 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2209");
        end

       2210 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2210");
        end

       2211 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2211");
        end

       2212 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2212");
        end

       2213 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2213");
        end

       2214 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2214");
        end

       2215 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2215");
        end

       2216 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2216");
        end

       2217 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2217");
        end

       2218 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2218");
        end

       2219 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2219");
        end

       2220 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2220");
        end

       2221 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2221");
        end

       2222 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2222");
        end

       2223 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2223");
        end

       2224 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2224");
        end

       2225 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2225");
        end

       2226 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2226");
        end

       2227 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2227");
        end

       2228 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2228");
        end

       2229 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2229");
        end

       2230 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2230");
        end

       2231 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2231");
        end

       2232 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2232");
        end

       2233 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2233");
        end

       2234 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2234");
        end

       2235 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2235");
        end

       2236 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2236");
        end

       2237 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2237");
        end

       2238 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2238");
        end

       2239 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2239");
        end

       2240 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2240");
        end

       2241 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2241");
        end

       2242 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2242");
        end

       2243 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2243");
        end

       2244 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2244");
        end

       2245 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2245");
        end

       2246 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2246");
        end

       2247 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2247");
        end

       2248 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2248");
        end

       2249 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2249");
        end

       2250 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2250");
        end

       2251 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2251");
        end

       2252 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2252");
        end

       2253 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2253");
        end

       2254 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2254");
        end

       2255 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2255");
        end

       2256 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2256");
        end

       2257 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2257");
        end

       2258 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2258");
        end

       2259 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2259");
        end

       2260 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2260");
        end

       2261 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2261");
        end

       2262 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2262");
        end

       2263 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2263");
        end

       2264 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2264");
        end

       2265 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2265");
        end

       2266 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2266");
        end

       2267 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2267");
        end

       2268 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2268");
        end

       2269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2269");
        end

       2270 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2270");
        end

       2271 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2271");
        end

       2272 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2272");
        end

       2273 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2273");
        end

       2274 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2274");
        end

       2275 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2275");
        end

       2276 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2276");
        end

       2277 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2277");
        end

       2278 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2278");
        end

       2279 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2279");
        end

       2280 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2280");
        end

       2281 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2281");
        end

       2282 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2282");
        end

       2283 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2283");
        end

       2284 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2284");
        end

       2285 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2285");
        end

       2286 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2286");
        end

       2287 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2287");
        end

       2288 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2288");
        end

       2289 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2289");
        end

       2290 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2290");
        end

       2291 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2291");
        end

       2292 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2292");
        end

       2293 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2293");
        end

       2294 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2294");
        end

       2295 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2295");
        end

       2296 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2296");
        end

       2297 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2297");
        end

       2298 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2298");
        end

       2299 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2299");
        end

       2300 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2300");
        end

       2301 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2301");
        end

       2302 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2302");
        end

       2303 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2303");
        end

       2304 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2304");
        end

       2305 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2305");
        end

       2306 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2306");
        end

       2307 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2307");
        end

       2308 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2308");
        end

       2309 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2309");
        end

       2310 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2310");
        end

       2311 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2311");
        end

       2312 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2312");
        end

       2313 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2313");
        end

       2314 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2314");
        end

       2315 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2315");
        end

       2316 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2317;
        end

       2317 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[142] = 1;
              ip = 2318;
        end

       2318 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2321;
        end

       2319 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2320;
        end

       2320 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[142] = 0;
              ip = 2321;
        end

       2321 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2322;
        end

       2322 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[142] != 0 ? 2324 : 2323;
        end

       2323 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[26] = localMem[141];
              ip = 2324;
        end

       2324 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2325;
        end

       2325 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3370;
        end

       2326 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2326");
        end

       2327 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2327");
        end

       2328 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2328");
        end

       2329 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2329");
        end

       2330 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2330");
        end

       2331 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2331");
        end

       2332 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2332");
        end

       2333 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2333");
        end

       2334 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  2334");
        end

       2335 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2335");
        end

       2336 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2336");
        end

       2337 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2337");
        end

       2338 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2338");
        end

       2339 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  2339");
        end

       2340 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2340");
        end

       2341 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2341");
        end

       2342 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2342");
        end

       2343 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2343");
        end

       2344 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2344");
        end

       2345 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2345");
        end

       2346 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2346");
        end

       2347 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2347");
        end

       2348 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  2348");
        end

       2349 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2349");
        end

       2350 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2350");
        end

       2351 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2351");
        end

       2352 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2352");
        end

       2353 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2353");
        end

       2354 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2354");
        end

       2355 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed  2355");
        end

       2356 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2356");
        end

       2357 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2357");
        end

       2358 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2358");
        end

       2359 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2359");
        end

       2360 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2360");
        end

       2361 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2361");
        end

       2362 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2362");
        end

       2363 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2363");
        end

       2364 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2364");
        end

       2365 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  2365");
        end

       2366 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  2366");
        end

       2367 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2367");
        end

       2368 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2368");
        end

       2369 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2369");
        end

       2370 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2370");
        end

       2371 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2371");
        end

       2372 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2372");
        end

       2373 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2373");
        end

       2374 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2374");
        end

       2375 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2375");
        end

       2376 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2376");
        end

       2377 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2377");
        end

       2378 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2378");
        end

       2379 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2379");
        end

       2380 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2380");
        end

       2381 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2381");
        end

       2382 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2382");
        end

       2383 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2383");
        end

       2384 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2384");
        end

       2385 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2385");
        end

       2386 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2386");
        end

       2387 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2387");
        end

       2388 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2388");
        end

       2389 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2389");
        end

       2390 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2390");
        end

       2391 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2391");
        end

       2392 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2392");
        end

       2393 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2393");
        end

       2394 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2394");
        end

       2395 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2395");
        end

       2396 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2396");
        end

       2397 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2397");
        end

       2398 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2398");
        end

       2399 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2399");
        end

       2400 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2400");
        end

       2401 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2401");
        end

       2402 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2402");
        end

       2403 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2403");
        end

       2404 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2404");
        end

       2405 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2405");
        end

       2406 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2406");
        end

       2407 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2407");
        end

       2408 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2408");
        end

       2409 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2409");
        end

       2410 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2410");
        end

       2411 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2411");
        end

       2412 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
          // $display("Should not be executed  2412");
        end

       2413 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2413");
        end

       2414 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
          // $display("Should not be executed  2414");
        end

       2415 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2415");
        end

       2416 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2416");
        end

       2417 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2417");
        end

       2418 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2418");
        end

       2419 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2419");
        end

       2420 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2420");
        end

       2421 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2421");
        end

       2422 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  2422");
        end

       2423 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2423");
        end

       2424 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2424");
        end

       2425 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2425");
        end

       2426 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2426");
        end

       2427 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2427");
        end

       2428 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2428");
        end

       2429 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2429");
        end

       2430 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2430");
        end

       2431 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2431");
        end

       2432 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2432");
        end

       2433 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2433");
        end

       2434 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2434");
        end

       2435 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2435");
        end

       2436 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2436");
        end

       2437 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2437");
        end

       2438 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2438");
        end

       2439 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2439");
        end

       2440 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2440");
        end

       2441 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2441");
        end

       2442 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2442");
        end

       2443 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2443");
        end

       2444 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2444");
        end

       2445 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2445");
        end

       2446 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2446");
        end

       2447 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2447");
        end

       2448 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2448");
        end

       2449 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2449");
        end

       2450 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2450");
        end

       2451 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2451");
        end

       2452 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2452");
        end

       2453 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2453");
        end

       2454 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2454");
        end

       2455 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2455");
        end

       2456 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2456");
        end

       2457 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2457");
        end

       2458 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2458");
        end

       2459 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2459");
        end

       2460 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2460");
        end

       2461 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2461");
        end

       2462 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2462");
        end

       2463 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2463");
        end

       2464 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2464");
        end

       2465 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2465");
        end

       2466 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2466");
        end

       2467 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2467");
        end

       2468 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2468");
        end

       2469 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2469");
        end

       2470 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2470");
        end

       2471 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2471");
        end

       2472 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2472");
        end

       2473 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2473");
        end

       2474 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2474");
        end

       2475 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2475");
        end

       2476 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2476");
        end

       2477 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2477");
        end

       2478 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2478");
        end

       2479 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2479");
        end

       2480 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2480");
        end

       2481 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2481");
        end

       2482 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2482");
        end

       2483 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2483");
        end

       2484 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2484");
        end

       2485 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2485");
        end

       2486 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2486");
        end

       2487 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2487");
        end

       2488 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  2488");
        end

       2489 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  2489");
        end

       2490 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2490");
        end

       2491 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2491");
        end

       2492 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2492");
        end

       2493 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2493");
        end

       2494 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2494");
        end

       2495 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2495");
        end

       2496 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2496");
        end

       2497 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2497");
        end

       2498 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2498");
        end

       2499 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2499");
        end

       2500 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2500");
        end

       2501 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2501");
        end

       2502 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2502");
        end

       2503 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2503");
        end

       2504 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2504");
        end

       2505 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2505");
        end

       2506 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2506");
        end

       2507 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2507");
        end

       2508 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2508");
        end

       2509 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2509");
        end

       2510 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2510");
        end

       2511 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2511");
        end

       2512 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2512");
        end

       2513 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2513");
        end

       2514 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2514");
        end

       2515 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2515");
        end

       2516 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2516");
        end

       2517 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2517");
        end

       2518 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2518");
        end

       2519 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2519");
        end

       2520 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2520");
        end

       2521 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2521");
        end

       2522 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2522");
        end

       2523 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2523");
        end

       2524 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2524");
        end

       2525 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2525");
        end

       2526 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2526");
        end

       2527 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2527");
        end

       2528 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2528");
        end

       2529 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2529");
        end

       2530 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2530");
        end

       2531 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2531");
        end

       2532 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2532");
        end

       2533 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2533");
        end

       2534 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2534");
        end

       2535 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2535");
        end

       2536 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2536");
        end

       2537 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2537");
        end

       2538 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2538");
        end

       2539 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2539");
        end

       2540 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2540");
        end

       2541 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2541");
        end

       2542 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2542");
        end

       2543 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2543");
        end

       2544 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2544");
        end

       2545 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2545");
        end

       2546 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2546");
        end

       2547 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2547");
        end

       2548 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2548");
        end

       2549 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2549");
        end

       2550 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2550");
        end

       2551 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2551");
        end

       2552 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2552");
        end

       2553 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2553");
        end

       2554 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2554");
        end

       2555 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2555");
        end

       2556 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2556");
        end

       2557 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2557");
        end

       2558 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2558");
        end

       2559 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2559");
        end

       2560 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2560");
        end

       2561 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2561");
        end

       2562 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2562");
        end

       2563 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2563");
        end

       2564 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2564");
        end

       2565 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2565");
        end

       2566 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2566");
        end

       2567 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2567");
        end

       2568 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2568");
        end

       2569 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2569");
        end

       2570 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2570");
        end

       2571 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2571");
        end

       2572 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2572");
        end

       2573 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2573");
        end

       2574 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2574");
        end

       2575 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2575");
        end

       2576 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2576");
        end

       2577 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2577");
        end

       2578 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2578");
        end

       2579 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2579");
        end

       2580 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2580");
        end

       2581 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2581");
        end

       2582 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2582");
        end

       2583 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2583");
        end

       2584 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2584");
        end

       2585 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2585");
        end

       2586 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2586");
        end

       2587 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2587");
        end

       2588 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2588");
        end

       2589 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2589");
        end

       2590 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2590");
        end

       2591 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2591");
        end

       2592 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2592");
        end

       2593 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2593");
        end

       2594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2594");
        end

       2595 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2595");
        end

       2596 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2596");
        end

       2597 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2597");
        end

       2598 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2598");
        end

       2599 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2599");
        end

       2600 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2600");
        end

       2601 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2601");
        end

       2602 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2602");
        end

       2603 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2603");
        end

       2604 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2604");
        end

       2605 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2605");
        end

       2606 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2606");
        end

       2607 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2607");
        end

       2608 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2608");
        end

       2609 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2609");
        end

       2610 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2610");
        end

       2611 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2611");
        end

       2612 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2612");
        end

       2613 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2613");
        end

       2614 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2614");
        end

       2615 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2615");
        end

       2616 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2616");
        end

       2617 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2617");
        end

       2618 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2618");
        end

       2619 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2619");
        end

       2620 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2620");
        end

       2621 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2621");
        end

       2622 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2622");
        end

       2623 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2623");
        end

       2624 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2624");
        end

       2625 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2625");
        end

       2626 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2626");
        end

       2627 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2627");
        end

       2628 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2628");
        end

       2629 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2629");
        end

       2630 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2630");
        end

       2631 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2631");
        end

       2632 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2632");
        end

       2633 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2633");
        end

       2634 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2634");
        end

       2635 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2635");
        end

       2636 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2636");
        end

       2637 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2637");
        end

       2638 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2638");
        end

       2639 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2639");
        end

       2640 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2640");
        end

       2641 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2641");
        end

       2642 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2642");
        end

       2643 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2643");
        end

       2644 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2644");
        end

       2645 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2645");
        end

       2646 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2646");
        end

       2647 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2647");
        end

       2648 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2648");
        end

       2649 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2649");
        end

       2650 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2650");
        end

       2651 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2651");
        end

       2652 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2652");
        end

       2653 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2653");
        end

       2654 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2654");
        end

       2655 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2655");
        end

       2656 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2656");
        end

       2657 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2657");
        end

       2658 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2658");
        end

       2659 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2659");
        end

       2660 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2660");
        end

       2661 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2661");
        end

       2662 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2662");
        end

       2663 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2663");
        end

       2664 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2664");
        end

       2665 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  2665");
        end

       2666 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2666");
        end

       2667 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2667");
        end

       2668 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2668");
        end

       2669 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2669");
        end

       2670 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2670");
        end

       2671 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2671");
        end

       2672 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2672");
        end

       2673 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2673");
        end

       2674 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2674");
        end

       2675 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2675");
        end

       2676 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2676");
        end

       2677 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2677");
        end

       2678 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2678");
        end

       2679 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2679");
        end

       2680 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2680");
        end

       2681 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2681");
        end

       2682 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2682");
        end

       2683 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2683");
        end

       2684 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2684");
        end

       2685 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2685");
        end

       2686 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2686");
        end

       2687 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2687");
        end

       2688 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2688");
        end

       2689 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2689");
        end

       2690 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2690");
        end

       2691 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2691");
        end

       2692 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2692");
        end

       2693 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2693");
        end

       2694 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2694");
        end

       2695 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2695");
        end

       2696 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2696");
        end

       2697 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2697");
        end

       2698 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2698");
        end

       2699 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2699");
        end

       2700 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2700");
        end

       2701 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2701");
        end

       2702 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2702");
        end

       2703 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2703");
        end

       2704 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2704");
        end

       2705 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2705");
        end

       2706 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2706");
        end

       2707 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2707");
        end

       2708 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2708");
        end

       2709 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2709");
        end

       2710 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2710");
        end

       2711 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2711");
        end

       2712 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2712");
        end

       2713 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2713");
        end

       2714 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2714");
        end

       2715 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2715");
        end

       2716 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2716");
        end

       2717 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2717");
        end

       2718 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2718");
        end

       2719 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2719");
        end

       2720 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2720");
        end

       2721 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2721");
        end

       2722 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2722");
        end

       2723 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2723");
        end

       2724 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2724");
        end

       2725 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2725");
        end

       2726 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2726");
        end

       2727 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2727");
        end

       2728 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2728");
        end

       2729 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2729");
        end

       2730 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2730");
        end

       2731 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2731");
        end

       2732 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2732");
        end

       2733 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2733");
        end

       2734 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2734");
        end

       2735 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2735");
        end

       2736 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2736");
        end

       2737 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2737");
        end

       2738 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2738");
        end

       2739 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2739");
        end

       2740 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2740");
        end

       2741 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2741");
        end

       2742 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2742");
        end

       2743 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2743");
        end

       2744 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2744");
        end

       2745 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2745");
        end

       2746 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  2746");
        end

       2747 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2747");
        end

       2748 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2748");
        end

       2749 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2749");
        end

       2750 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2750");
        end

       2751 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2751");
        end

       2752 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2752");
        end

       2753 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2753");
        end

       2754 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  2754");
        end

       2755 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2755");
        end

       2756 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2756");
        end

       2757 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2757");
        end

       2758 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2758");
        end

       2759 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  2759");
        end

       2760 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2760");
        end

       2761 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2761");
        end

       2762 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2762");
        end

       2763 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2763");
        end

       2764 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2764");
        end

       2765 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2765");
        end

       2766 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2766");
        end

       2767 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2767");
        end

       2768 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2768");
        end

       2769 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2769");
        end

       2770 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2770");
        end

       2771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2771");
        end

       2772 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2772");
        end

       2773 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2773");
        end

       2774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2774");
        end

       2775 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2775");
        end

       2776 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2776");
        end

       2777 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2777");
        end

       2778 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2778");
        end

       2779 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2779");
        end

       2780 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2780");
        end

       2781 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2781");
        end

       2782 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2782");
        end

       2783 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2783");
        end

       2784 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2784");
        end

       2785 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2785");
        end

       2786 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2786");
        end

       2787 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2787");
        end

       2788 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2788");
        end

       2789 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2789");
        end

       2790 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2790");
        end

       2791 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2791");
        end

       2792 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2792");
        end

       2793 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2793");
        end

       2794 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2794");
        end

       2795 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2795");
        end

       2796 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2796");
        end

       2797 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2797");
        end

       2798 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2798");
        end

       2799 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2799");
        end

       2800 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2800");
        end

       2801 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2801");
        end

       2802 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2802");
        end

       2803 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2803");
        end

       2804 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2804");
        end

       2805 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2805");
        end

       2806 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2806");
        end

       2807 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2807");
        end

       2808 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2808");
        end

       2809 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2809");
        end

       2810 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2810");
        end

       2811 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2811");
        end

       2812 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2812");
        end

       2813 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2813");
        end

       2814 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2814");
        end

       2815 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2815");
        end

       2816 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2816");
        end

       2817 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2817");
        end

       2818 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2818");
        end

       2819 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2819");
        end

       2820 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2820");
        end

       2821 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2821");
        end

       2822 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2822");
        end

       2823 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2823");
        end

       2824 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2824");
        end

       2825 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2825");
        end

       2826 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2826");
        end

       2827 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2827");
        end

       2828 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2828");
        end

       2829 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2829");
        end

       2830 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2830");
        end

       2831 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2831");
        end

       2832 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2832");
        end

       2833 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2833");
        end

       2834 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2834");
        end

       2835 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2835");
        end

       2836 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2836");
        end

       2837 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2837");
        end

       2838 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2838");
        end

       2839 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2839");
        end

       2840 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2840");
        end

       2841 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2841");
        end

       2842 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2842");
        end

       2843 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2843");
        end

       2844 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2844");
        end

       2845 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2845");
        end

       2846 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2846");
        end

       2847 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2847");
        end

       2848 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2848");
        end

       2849 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2849");
        end

       2850 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2850");
        end

       2851 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2851");
        end

       2852 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2852");
        end

       2853 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2853");
        end

       2854 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2854");
        end

       2855 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2855");
        end

       2856 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2856");
        end

       2857 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2857");
        end

       2858 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2858");
        end

       2859 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2859");
        end

       2860 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2860");
        end

       2861 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2861");
        end

       2862 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2862");
        end

       2863 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2863");
        end

       2864 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2864");
        end

       2865 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2865");
        end

       2866 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2866");
        end

       2867 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2867");
        end

       2868 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2868");
        end

       2869 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2869");
        end

       2870 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2870");
        end

       2871 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2871");
        end

       2872 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2872");
        end

       2873 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2873");
        end

       2874 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2874");
        end

       2875 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2875");
        end

       2876 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2876");
        end

       2877 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2877");
        end

       2878 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2878");
        end

       2879 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2879");
        end

       2880 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2880");
        end

       2881 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2881");
        end

       2882 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2882");
        end

       2883 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2883");
        end

       2884 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2884");
        end

       2885 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2885");
        end

       2886 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2886");
        end

       2887 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2887");
        end

       2888 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2888");
        end

       2889 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2889");
        end

       2890 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2890");
        end

       2891 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2891");
        end

       2892 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2892");
        end

       2893 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2893");
        end

       2894 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2894");
        end

       2895 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2895");
        end

       2896 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2896");
        end

       2897 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2897");
        end

       2898 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2898");
        end

       2899 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2899");
        end

       2900 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2900");
        end

       2901 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2901");
        end

       2902 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2902");
        end

       2903 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2903");
        end

       2904 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2904");
        end

       2905 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2905");
        end

       2906 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2906");
        end

       2907 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2907");
        end

       2908 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2908");
        end

       2909 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2909");
        end

       2910 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2910");
        end

       2911 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2911");
        end

       2912 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2912");
        end

       2913 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2913");
        end

       2914 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2914");
        end

       2915 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2915");
        end

       2916 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2916");
        end

       2917 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2917");
        end

       2918 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2918");
        end

       2919 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2919");
        end

       2920 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2920");
        end

       2921 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2921");
        end

       2922 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2922");
        end

       2923 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2923");
        end

       2924 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2924");
        end

       2925 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2925");
        end

       2926 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2926");
        end

       2927 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2927");
        end

       2928 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2928");
        end

       2929 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2929");
        end

       2930 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2930");
        end

       2931 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2931");
        end

       2932 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2932");
        end

       2933 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2933");
        end

       2934 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2934");
        end

       2935 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2935");
        end

       2936 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2936");
        end

       2937 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2937");
        end

       2938 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2938");
        end

       2939 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2939");
        end

       2940 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2940");
        end

       2941 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2941");
        end

       2942 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2942");
        end

       2943 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2943");
        end

       2944 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2944");
        end

       2945 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2945");
        end

       2946 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2946");
        end

       2947 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2947");
        end

       2948 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2948");
        end

       2949 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2949");
        end

       2950 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2950");
        end

       2951 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2951");
        end

       2952 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2952");
        end

       2953 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2953");
        end

       2954 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2954");
        end

       2955 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2955");
        end

       2956 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2956");
        end

       2957 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2957");
        end

       2958 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2958");
        end

       2959 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2959");
        end

       2960 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2960");
        end

       2961 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2961");
        end

       2962 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2962");
        end

       2963 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2963");
        end

       2964 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2964");
        end

       2965 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2965");
        end

       2966 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2966");
        end

       2967 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  2967");
        end

       2968 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  2968");
        end

       2969 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2969");
        end

       2970 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2970");
        end

       2971 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2971");
        end

       2972 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2972");
        end

       2973 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2973");
        end

       2974 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2974");
        end

       2975 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2975");
        end

       2976 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2976");
        end

       2977 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2977");
        end

       2978 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2978");
        end

       2979 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2979");
        end

       2980 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2980");
        end

       2981 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2981");
        end

       2982 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2982");
        end

       2983 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2983");
        end

       2984 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2984");
        end

       2985 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2985");
        end

       2986 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2986");
        end

       2987 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2987");
        end

       2988 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2988");
        end

       2989 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2989");
        end

       2990 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2990");
        end

       2991 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2991");
        end

       2992 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2992");
        end

       2993 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2993");
        end

       2994 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2994");
        end

       2995 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2995");
        end

       2996 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2996");
        end

       2997 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2997");
        end

       2998 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2998");
        end

       2999 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2999");
        end

       3000 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3000");
        end

       3001 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3001");
        end

       3002 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3002");
        end

       3003 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3003");
        end

       3004 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3004");
        end

       3005 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3005");
        end

       3006 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3006");
        end

       3007 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3007");
        end

       3008 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3008");
        end

       3009 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3009");
        end

       3010 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3010");
        end

       3011 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3011");
        end

       3012 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3012");
        end

       3013 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3013");
        end

       3014 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3014");
        end

       3015 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3015");
        end

       3016 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3016");
        end

       3017 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3017");
        end

       3018 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3018");
        end

       3019 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3019");
        end

       3020 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3020");
        end

       3021 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3021");
        end

       3022 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3022");
        end

       3023 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3023");
        end

       3024 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3024");
        end

       3025 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3025");
        end

       3026 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3026");
        end

       3027 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3027");
        end

       3028 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3028");
        end

       3029 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3029");
        end

       3030 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3030");
        end

       3031 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3031");
        end

       3032 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3032");
        end

       3033 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3033");
        end

       3034 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3034");
        end

       3035 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3035");
        end

       3036 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3036");
        end

       3037 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3037");
        end

       3038 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3038");
        end

       3039 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3039");
        end

       3040 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3040");
        end

       3041 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3041");
        end

       3042 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3042");
        end

       3043 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3043");
        end

       3044 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3044");
        end

       3045 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3045");
        end

       3046 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3046");
        end

       3047 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3047");
        end

       3048 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3048");
        end

       3049 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3049");
        end

       3050 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3050");
        end

       3051 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3051");
        end

       3052 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3052");
        end

       3053 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3053");
        end

       3054 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3054");
        end

       3055 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3055");
        end

       3056 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3056");
        end

       3057 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3057");
        end

       3058 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3058");
        end

       3059 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3059");
        end

       3060 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3060");
        end

       3061 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3061");
        end

       3062 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3062");
        end

       3063 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3063");
        end

       3064 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3064");
        end

       3065 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3065");
        end

       3066 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3066");
        end

       3067 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3067");
        end

       3068 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3068");
        end

       3069 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3069");
        end

       3070 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3070");
        end

       3071 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3071");
        end

       3072 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3072");
        end

       3073 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3073");
        end

       3074 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3074");
        end

       3075 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3075");
        end

       3076 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3076");
        end

       3077 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3077");
        end

       3078 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3078");
        end

       3079 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3079");
        end

       3080 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3080");
        end

       3081 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3081");
        end

       3082 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3082");
        end

       3083 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3083");
        end

       3084 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3084");
        end

       3085 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3085");
        end

       3086 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3086");
        end

       3087 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3087");
        end

       3088 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3088");
        end

       3089 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3089");
        end

       3090 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3090");
        end

       3091 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3091");
        end

       3092 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3092");
        end

       3093 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3093");
        end

       3094 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3094");
        end

       3095 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3095");
        end

       3096 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3096");
        end

       3097 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3097");
        end

       3098 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3098");
        end

       3099 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3099");
        end

       3100 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3100");
        end

       3101 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3101");
        end

       3102 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3102");
        end

       3103 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3103");
        end

       3104 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3104");
        end

       3105 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3105");
        end

       3106 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3106");
        end

       3107 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3107");
        end

       3108 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3108");
        end

       3109 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3109");
        end

       3110 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3110");
        end

       3111 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3111");
        end

       3112 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3112");
        end

       3113 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3113");
        end

       3114 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3114");
        end

       3115 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3115");
        end

       3116 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3116");
        end

       3117 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3117");
        end

       3118 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3118");
        end

       3119 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3119");
        end

       3120 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3120");
        end

       3121 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  3121");
        end

       3122 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3122");
        end

       3123 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3123");
        end

       3124 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3124");
        end

       3125 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3125");
        end

       3126 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3126");
        end

       3127 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3127");
        end

       3128 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3128");
        end

       3129 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3129");
        end

       3130 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3130");
        end

       3131 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3131");
        end

       3132 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3132");
        end

       3133 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3133");
        end

       3134 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3134");
        end

       3135 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3135");
        end

       3136 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3136");
        end

       3137 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3137");
        end

       3138 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3138");
        end

       3139 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3139");
        end

       3140 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3140");
        end

       3141 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3141");
        end

       3142 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3142");
        end

       3143 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3143");
        end

       3144 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3144");
        end

       3145 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3145");
        end

       3146 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3146");
        end

       3147 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3147");
        end

       3148 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3148");
        end

       3149 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3149");
        end

       3150 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3150");
        end

       3151 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3151");
        end

       3152 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  3152");
        end

       3153 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3153");
        end

       3154 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3154");
        end

       3155 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3155");
        end

       3156 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3156");
        end

       3157 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3157");
        end

       3158 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3158");
        end

       3159 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3159");
        end

       3160 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3160");
        end

       3161 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3161");
        end

       3162 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3162");
        end

       3163 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3163");
        end

       3164 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3164");
        end

       3165 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3165");
        end

       3166 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3166");
        end

       3167 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3167");
        end

       3168 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3168");
        end

       3169 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3169");
        end

       3170 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  3170");
        end

       3171 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3171");
        end

       3172 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3172");
        end

       3173 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3173");
        end

       3174 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3174");
        end

       3175 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3175");
        end

       3176 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3176");
        end

       3177 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3177");
        end

       3178 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3178");
        end

       3179 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3179");
        end

       3180 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3180");
        end

       3181 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3181");
        end

       3182 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3182");
        end

       3183 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3183");
        end

       3184 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3184");
        end

       3185 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3185");
        end

       3186 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3186");
        end

       3187 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3187");
        end

       3188 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3188");
        end

       3189 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3189");
        end

       3190 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3190");
        end

       3191 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3191");
        end

       3192 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3192");
        end

       3193 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3193");
        end

       3194 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3194");
        end

       3195 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3195");
        end

       3196 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3196");
        end

       3197 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3197");
        end

       3198 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3198");
        end

       3199 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3199");
        end

       3200 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3200");
        end

       3201 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3201");
        end

       3202 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3202");
        end

       3203 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3203");
        end

       3204 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3204");
        end

       3205 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3205");
        end

       3206 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3206");
        end

       3207 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3207");
        end

       3208 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3208");
        end

       3209 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3209");
        end

       3210 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3210");
        end

       3211 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3211");
        end

       3212 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3212");
        end

       3213 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3213");
        end

       3214 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3214");
        end

       3215 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3215");
        end

       3216 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3216");
        end

       3217 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3217");
        end

       3218 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3218");
        end

       3219 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3219");
        end

       3220 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3220");
        end

       3221 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3221");
        end

       3222 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3222");
        end

       3223 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3223");
        end

       3224 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3224");
        end

       3225 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3225");
        end

       3226 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3226");
        end

       3227 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3227");
        end

       3228 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3228");
        end

       3229 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3229");
        end

       3230 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3230");
        end

       3231 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3231");
        end

       3232 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3232");
        end

       3233 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3233");
        end

       3234 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3234");
        end

       3235 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3235");
        end

       3236 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3236");
        end

       3237 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3237");
        end

       3238 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3238");
        end

       3239 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3239");
        end

       3240 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3240");
        end

       3241 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3241");
        end

       3242 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3242");
        end

       3243 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3243");
        end

       3244 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3244");
        end

       3245 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3245");
        end

       3246 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3246");
        end

       3247 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3247");
        end

       3248 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3248");
        end

       3249 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3249");
        end

       3250 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3250");
        end

       3251 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3251");
        end

       3252 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3252");
        end

       3253 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3253");
        end

       3254 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3254");
        end

       3255 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3255");
        end

       3256 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3256");
        end

       3257 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3257");
        end

       3258 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3258");
        end

       3259 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3259");
        end

       3260 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3260");
        end

       3261 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3261");
        end

       3262 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3262");
        end

       3263 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3263");
        end

       3264 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3264");
        end

       3265 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3265");
        end

       3266 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3266");
        end

       3267 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3267");
        end

       3268 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3268");
        end

       3269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3269");
        end

       3270 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3270");
        end

       3271 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3271");
        end

       3272 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3272");
        end

       3273 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3273");
        end

       3274 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3274");
        end

       3275 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3275");
        end

       3276 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3276");
        end

       3277 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3277");
        end

       3278 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3278");
        end

       3279 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3279");
        end

       3280 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3280");
        end

       3281 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3281");
        end

       3282 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3282");
        end

       3283 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3283");
        end

       3284 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3284");
        end

       3285 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3285");
        end

       3286 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3286");
        end

       3287 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3287");
        end

       3288 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3288");
        end

       3289 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3289");
        end

       3290 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3290");
        end

       3291 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3291");
        end

       3292 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3292");
        end

       3293 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3293");
        end

       3294 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3294");
        end

       3295 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3295");
        end

       3296 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3296");
        end

       3297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3297");
        end

       3298 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3298");
        end

       3299 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3299");
        end

       3300 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3300");
        end

       3301 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3301");
        end

       3302 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3302");
        end

       3303 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3303");
        end

       3304 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3304");
        end

       3305 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3305");
        end

       3306 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3306");
        end

       3307 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3307");
        end

       3308 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3308");
        end

       3309 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3309");
        end

       3310 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3310");
        end

       3311 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3311");
        end

       3312 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3312");
        end

       3313 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3313");
        end

       3314 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3314");
        end

       3315 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3315");
        end

       3316 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3316");
        end

       3317 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3317");
        end

       3318 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3318");
        end

       3319 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3319");
        end

       3320 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3320");
        end

       3321 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3321");
        end

       3322 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3322");
        end

       3323 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3323");
        end

       3324 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3324");
        end

       3325 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3325");
        end

       3326 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3326");
        end

       3327 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3327");
        end

       3328 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3328");
        end

       3329 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3329");
        end

       3330 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3330");
        end

       3331 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3331");
        end

       3332 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3332");
        end

       3333 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3333");
        end

       3334 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3334");
        end

       3335 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3335");
        end

       3336 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3336");
        end

       3337 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3337");
        end

       3338 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3338");
        end

       3339 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3339");
        end

       3340 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3340");
        end

       3341 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3341");
        end

       3342 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3342");
        end

       3343 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3343");
        end

       3344 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3344");
        end

       3345 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3345");
        end

       3346 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3346");
        end

       3347 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3347");
        end

       3348 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3348");
        end

       3349 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3349");
        end

       3350 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3350");
        end

       3351 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3351");
        end

       3352 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3352");
        end

       3353 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3353");
        end

       3354 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3354");
        end

       3355 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3355");
        end

       3356 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3356");
        end

       3357 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3357");
        end

       3358 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3358");
        end

       3359 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3359");
        end

       3360 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3360");
        end

       3361 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3361");
        end

       3362 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3362");
        end

       3363 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3363");
        end

       3364 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3364");
        end

       3365 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3365");
        end

       3366 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3366");
        end

       3367 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  3367");
        end

       3368 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3368");
        end

       3369 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3369");
        end

       3370 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3371;
        end

       3371 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[134] = localMem[134] + 1;
              ip = 3372;
        end

       3372 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1293;
        end

       3373 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3373");
        end

       3374 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  3374");
        end

       3375 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3375");
        end

       3376 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3376");
        end

       3377 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3378;
        end

       3378 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3379;
        end

       3379 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3380;
              heapClock = 1;
        end

       3380 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3381;
        end

       3381 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[970] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3382;
              heapClock = 1;
        end

       3382 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3383;
        end

       3383 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[362] = localMem[970];
              ip = 3384;
        end

       3384 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3385;
        end

       3385 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3386;
              heapClock = 1;
        end

       3386 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3387;
        end

       3387 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[971] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3388;
              heapClock = 1;
        end

       3388 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3389;
        end

       3389 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[363] = localMem[971];
              ip = 3390;
        end

       3390 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3391;
        end

       3391 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3392;
              heapClock = 1;
        end

       3392 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3393;
        end

       3393 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[972] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3394;
              heapClock = 1;
        end

       3394 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3395;
        end

       3395 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[364] = localMem[972];
              ip = 3396;
        end

       3396 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[363] != 1 ? 3408 : 3397;
        end

       3397 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3397");
        end

       3398 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3398");
        end

       3399 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3399");
        end

       3400 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3400");
        end

       3401 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3401");
        end

       3402 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3402");
        end

       3403 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3403");
        end

       3404 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3404");
        end

       3405 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3405");
        end

       3406 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3406");
        end

       3407 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3407");
        end

       3408 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3409;
        end

       3409 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[363] != 2 ? 3439 : 3410;
        end

       3410 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[366] = localMem[364] + 1;
              ip = 3411;
        end

       3411 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3412;
        end

       3412 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3413;
              heapClock = 1;
        end

       3413 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3414;
        end

       3414 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[975] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3415;
              heapClock = 1;
        end

       3415 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3416;
        end

       3416 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[367] = localMem[975];
              ip = 3417;
        end

       3417 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3418;
        end

       3418 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[1];
              heapArray  = localMem[367];
              heapIndex  = localMem[366];
              ip = 3419;
              heapClock = 1;
        end

       3419 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3420;
        end

       3420 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3421;
        end

       3421 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3422;
              heapClock = 1;
        end

       3422 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3423;
        end

       3423 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[976] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3424;
              heapClock = 1;
        end

       3424 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3425;
        end

       3425 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[368] = localMem[976];
              ip = 3426;
        end

       3426 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3427;
        end

       3427 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[2];
              heapArray  = localMem[368];
              heapIndex  = localMem[366];
              ip = 3428;
              heapClock = 1;
        end

       3428 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3429;
        end

       3429 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3430;
        end

       3430 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3431;
              heapClock = 1;
        end

       3431 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3432;
        end

       3432 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[977] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3433;
              heapClock = 1;
        end

       3433 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3434;
        end

       3434 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[978] = localMem[977] + 1;
              ip = 3435;
        end

       3435 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3436;
        end

       3436 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[362];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[978];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3437;
              heapClock = 1;
        end

       3437 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3438;
        end

       3438 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3467;
        end

       3439 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3439");
        end

       3440 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3440");
        end

       3441 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3441");
        end

       3442 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3442");
        end

       3443 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3443");
        end

       3444 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3444");
        end

       3445 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3445");
        end

       3446 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3446");
        end

       3447 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  3447");
        end

       3448 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3448");
        end

       3449 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3449");
        end

       3450 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3450");
        end

       3451 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3451");
        end

       3452 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3452");
        end

       3453 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3453");
        end

       3454 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3454");
        end

       3455 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3455");
        end

       3456 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  3456");
        end

       3457 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3457");
        end

       3458 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3458");
        end

       3459 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3459");
        end

       3460 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3460");
        end

       3461 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3461");
        end

       3462 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3462");
        end

       3463 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3463");
        end

       3464 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3464");
        end

       3465 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3465");
        end

       3466 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3466");
        end

       3467 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3468;
        end

       3468 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3469;
        end

       3469 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3470;
              heapClock = 1;
        end

       3470 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3471;
        end

       3471 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[983] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3472;
              heapClock = 1;
        end

       3472 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3473;
        end

       3473 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[984] = localMem[983] + 1;
              ip = 3474;
        end

       3474 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3475;
        end

       3475 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[984];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3476;
              heapClock = 1;
        end

       3476 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3477;
        end

       3477 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3478;
        end

       3478 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3479;
        end

       3479 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3480;
              heapClock = 1;
        end

       3480 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3481;
        end

       3481 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[985] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3482;
              heapClock = 1;
        end

       3482 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3483;
        end

       3483 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[372] = localMem[985];
              ip = 3484;
        end

       3484 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3485;
        end

       3485 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3486;
              heapClock = 1;
        end

       3486 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3487;
        end

       3487 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[986] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3488;
              heapClock = 1;
        end

       3488 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3489;
        end

       3489 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[373] = localMem[986];
              ip = 3490;
        end

       3490 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3491;
        end

       3491 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3492;
              heapClock = 1;
        end

       3492 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3493;
        end

       3493 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[987] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3494;
              heapClock = 1;
        end

       3494 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3495;
        end

       3495 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[374] = localMem[987];
              ip = 3496;
        end

       3496 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[372] <  localMem[374] ? 4448 : 3497;
        end

       3497 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[375] = localMem[374];
              ip = 3498;
        end

       3498 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[375] = localMem[375] >> 1;
              ip = 3499;
              ip = 3499;
        end

       3499 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[376] = localMem[375] + 1;
              ip = 3500;
        end

       3500 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3501;
        end

       3501 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3502;
              heapClock = 1;
        end

       3502 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3503;
        end

       3503 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[988] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3504;
              heapClock = 1;
        end

       3504 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3505;
        end

       3505 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[377] = localMem[988];
              ip = 3506;
        end

       3506 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[377] == 0 ? 3925 : 3507;
        end

       3507 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3508;
        end

       3508 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3509;
              heapClock = 1;
        end

       3509 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3510;
        end

       3510 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[378] = heapOut;
              ip = 3511;
        end

       3511 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3512;
        end

       3512 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3513;
        end

       3513 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[989] = localMem[375];
              ip = 3514;
        end

       3514 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3515;
        end

       3515 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[989];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3516;
              heapClock = 1;
        end

       3516 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3517;
        end

       3517 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[990] = 0;
              ip = 3518;
        end

       3518 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3519;
        end

       3519 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[990];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3520;
              heapClock = 1;
        end

       3520 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3521;
        end

       3521 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3522;
        end

       3522 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3523;
              heapClock = 1;
        end

       3523 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3524;
        end

       3524 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[379] = heapOut;
              ip = 3525;
        end

       3525 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3526;
        end

       3526 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3527;
        end

       3527 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[991] = localMem[379];
              ip = 3528;
        end

       3528 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3529;
        end

       3529 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[991];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3530;
              heapClock = 1;
        end

       3530 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3531;
        end

       3531 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3532;
        end

       3532 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3533;
              heapClock = 1;
        end

       3533 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3534;
        end

       3534 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[380] = heapOut;
              ip = 3535;
        end

       3535 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3536;
        end

       3536 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3537;
        end

       3537 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[992] = localMem[380];
              ip = 3538;
        end

       3538 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3539;
        end

       3539 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[992];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3540;
              heapClock = 1;
        end

       3540 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3541;
        end

       3541 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[993] = 0;
              ip = 3542;
        end

       3542 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3543;
        end

       3543 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[993];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3544;
              heapClock = 1;
        end

       3544 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3545;
        end

       3545 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[994] = localMem[373];
              ip = 3546;
        end

       3546 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3547;
        end

       3547 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[994];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3548;
              heapClock = 1;
        end

       3548 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3549;
        end

       3549 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3550;
        end

       3550 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3551;
              heapClock = 1;
        end

       3551 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3552;
        end

       3552 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[995] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3553;
              heapClock = 1;
        end

       3553 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3554;
        end

       3554 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[996] = localMem[995] + 1;
              ip = 3555;
        end

       3555 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3556;
        end

       3556 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[373];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[996];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3557;
              heapClock = 1;
        end

       3557 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3558;
        end

       3558 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3559;
        end

       3559 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3560;
              heapClock = 1;
        end

       3560 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3561;
        end

       3561 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[997] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3562;
              heapClock = 1;
        end

       3562 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3563;
        end

       3563 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[998] = localMem[997];
              ip = 3564;
        end

       3564 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3565;
        end

       3565 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[998];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3566;
              heapClock = 1;
        end

       3566 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3567;
        end

       3567 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3568;
        end

       3568 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3569;
              heapClock = 1;
        end

       3569 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3570;
        end

       3570 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[999] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3571;
              heapClock = 1;
        end

       3571 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3572;
        end

       3572 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[381] = !localMem[999];
              ip = 3573;
        end

       3573 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[381] != 0 ? 3683 : 3574;
        end

       3574 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3574");
        end

       3575 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  3575");
        end

       3576 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3576");
        end

       3577 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3577");
        end

       3578 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3578");
        end

       3579 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3579");
        end

       3580 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3580");
        end

       3581 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3581");
        end

       3582 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3582");
        end

       3583 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3583");
        end

       3584 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3584");
        end

       3585 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3585");
        end

       3586 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3586");
        end

       3587 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3587");
        end

       3588 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3588");
        end

       3589 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3589");
        end

       3590 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3590");
        end

       3591 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3591");
        end

       3592 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3592");
        end

       3593 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3593");
        end

       3594 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3594");
        end

       3595 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3595");
        end

       3596 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3596");
        end

       3597 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3597");
        end

       3598 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3598");
        end

       3599 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3599");
        end

       3600 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3600");
        end

       3601 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3601");
        end

       3602 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3602");
        end

       3603 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3603");
        end

       3604 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3604");
        end

       3605 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3605");
        end

       3606 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3606");
        end

       3607 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3607");
        end

       3608 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3608");
        end

       3609 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3609");
        end

       3610 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3610");
        end

       3611 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3611");
        end

       3612 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3612");
        end

       3613 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3613");
        end

       3614 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3614");
        end

       3615 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3615");
        end

       3616 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3616");
        end

       3617 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3617");
        end

       3618 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3618");
        end

       3619 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3619");
        end

       3620 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3620");
        end

       3621 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3621");
        end

       3622 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3622");
        end

       3623 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3623");
        end

       3624 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3624");
        end

       3625 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3625");
        end

       3626 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3626");
        end

       3627 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3627");
        end

       3628 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3628");
        end

       3629 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3629");
        end

       3630 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3630");
        end

       3631 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3631");
        end

       3632 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3632");
        end

       3633 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3633");
        end

       3634 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3634");
        end

       3635 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3635");
        end

       3636 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3636");
        end

       3637 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3637");
        end

       3638 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3638");
        end

       3639 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3639");
        end

       3640 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3640");
        end

       3641 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3641");
        end

       3642 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3642");
        end

       3643 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3643");
        end

       3644 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3644");
        end

       3645 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3645");
        end

       3646 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3646");
        end

       3647 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3647");
        end

       3648 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3648");
        end

       3649 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3649");
        end

       3650 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3650");
        end

       3651 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3651");
        end

       3652 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3652");
        end

       3653 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3653");
        end

       3654 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3654");
        end

       3655 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3655");
        end

       3656 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3656");
        end

       3657 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3657");
        end

       3658 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  3658");
        end

       3659 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3659");
        end

       3660 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3660");
        end

       3661 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3661");
        end

       3662 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3662");
        end

       3663 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3663");
        end

       3664 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3664");
        end

       3665 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3665");
        end

       3666 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3666");
        end

       3667 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3667");
        end

       3668 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3668");
        end

       3669 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3669");
        end

       3670 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3670");
        end

       3671 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3671");
        end

       3672 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3672");
        end

       3673 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3673");
        end

       3674 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3674");
        end

       3675 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3675");
        end

       3676 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3676");
        end

       3677 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3677");
        end

       3678 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3678");
        end

       3679 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3679");
        end

       3680 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3680");
        end

       3681 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3681");
        end

       3682 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3682");
        end

       3683 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3684;
        end

       3684 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3685;
        end

       3685 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3686;
              heapClock = 1;
        end

       3686 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3687;
        end

       3687 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1012] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3688;
              heapClock = 1;
        end

       3688 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3689;
        end

       3689 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[396] = localMem[1012];
              ip = 3690;
        end

       3690 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3691;
        end

       3691 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[378];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3692;
              heapClock = 1;
        end

       3692 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3693;
        end

       3693 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1013] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3694;
              heapClock = 1;
        end

       3694 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3695;
        end

       3695 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[397] = localMem[1013];
              ip = 3696;
        end

       3696 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3697;
        end

       3697 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3698;
        end

       3698 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[396];                                                 // Array to write to
              heapIndex  = localMem[376];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 3699;
              heapClock = 1;
        end

       3699 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3700;
        end

       3700 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[397];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[375];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 3701;
              heapClock = 1;
        end

       3701 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3702;
        end

       3702 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3703;
        end

       3703 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3704;
        end

       3704 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3705;
              heapClock = 1;
        end

       3705 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3706;
        end

       3706 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1014] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3707;
              heapClock = 1;
        end

       3707 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3708;
        end

       3708 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[398] = localMem[1014];
              ip = 3709;
        end

       3709 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3710;
        end

       3710 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[378];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3711;
              heapClock = 1;
        end

       3711 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3712;
        end

       3712 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1015] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3713;
              heapClock = 1;
        end

       3713 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3714;
        end

       3714 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[399] = localMem[1015];
              ip = 3715;
        end

       3715 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3716;
        end

       3716 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3717;
        end

       3717 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[398];                                                 // Array to write to
              heapIndex  = localMem[376];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 3718;
              heapClock = 1;
        end

       3718 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3719;
        end

       3719 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[399];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[375];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 3720;
              heapClock = 1;
        end

       3720 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3721;
        end

       3721 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3722;
        end

       3722 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3723;
        end

       3723 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1016] = localMem[375];
              ip = 3724;
        end

       3724 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3725;
        end

       3725 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[362];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1016];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3726;
              heapClock = 1;
        end

       3726 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3727;
        end

       3727 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1017] = localMem[377];
              ip = 3728;
        end

       3728 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3729;
        end

       3729 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1017];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3730;
              heapClock = 1;
        end

       3730 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3731;
        end

       3731 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3732;
        end

       3732 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3733;
              heapClock = 1;
        end

       3733 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3734;
        end

       3734 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1018] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3735;
              heapClock = 1;
        end

       3735 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3736;
        end

       3736 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[400] = localMem[1018];
              ip = 3737;
        end

       3737 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3738;
        end

       3738 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3739;
              heapClock = 1;
        end

       3739 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3740;
        end

       3740 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1019] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3741;
              heapClock = 1;
        end

       3741 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3742;
        end

       3742 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[401] = localMem[1019];
              ip = 3743;
        end

       3743 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3744;
        end

       3744 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[401];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[400];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3745;
              heapClock = 1;
        end

       3745 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3746;
        end

       3746 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1020] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3747;
              heapClock = 1;
        end

       3747 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3748;
        end

       3748 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[402] = localMem[1020];
              ip = 3749;
        end

       3749 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[402] != localMem[362] ? 3829 : 3750;
        end

       3750 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3751;
        end

       3751 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3752;
              heapClock = 1;
        end

       3752 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3753;
        end

       3753 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1021] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3754;
              heapClock = 1;
        end

       3754 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3755;
        end

       3755 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[403] = localMem[1021];
              ip = 3756;
        end

       3756 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3757;
        end

       3757 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[403];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[375];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3758;
              heapClock = 1;
        end

       3758 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3759;
        end

       3759 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1022] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3760;
              heapClock = 1;
        end

       3760 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3761;
        end

       3761 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[404] = localMem[1022];
              ip = 3762;
        end

       3762 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3763;
        end

       3763 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3764;
              heapClock = 1;
        end

       3764 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3765;
        end

       3765 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1023] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3766;
              heapClock = 1;
        end

       3766 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3767;
        end

       3767 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[405] = localMem[1023];
              ip = 3768;
        end

       3768 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1024] = localMem[404];
              ip = 3769;
        end

       3769 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3770;
        end

       3770 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[405];                                                // Array to write to
              heapIndex   = localMem[400];                                                // Index of element to write to
              heapIn      = localMem[1024];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3771;
              heapClock = 1;
        end

       3771 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3772;
        end

       3772 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3773;
        end

       3773 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3774;
              heapClock = 1;
        end

       3774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3775;
        end

       3775 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1025] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3776;
              heapClock = 1;
        end

       3776 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3777;
        end

       3777 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[406] = localMem[1025];
              ip = 3778;
        end

       3778 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3779;
        end

       3779 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[406];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[375];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3780;
              heapClock = 1;
        end

       3780 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3781;
        end

       3781 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1026] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3782;
              heapClock = 1;
        end

       3782 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3783;
        end

       3783 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[407] = localMem[1026];
              ip = 3784;
        end

       3784 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3785;
        end

       3785 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3786;
              heapClock = 1;
        end

       3786 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3787;
        end

       3787 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1027] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3788;
              heapClock = 1;
        end

       3788 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3789;
        end

       3789 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[408] = localMem[1027];
              ip = 3790;
        end

       3790 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1028] = localMem[407];
              ip = 3791;
        end

       3791 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3792;
        end

       3792 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[408];                                                // Array to write to
              heapIndex   = localMem[400];                                                // Index of element to write to
              heapIn      = localMem[1028];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3793;
              heapClock = 1;
        end

       3793 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3794;
        end

       3794 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3795;
        end

       3795 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3796;
              heapClock = 1;
        end

       3796 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3797;
        end

       3797 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1029] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3798;
              heapClock = 1;
        end

       3798 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3799;
        end

       3799 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[409] = localMem[1029];
              ip = 3800;
        end

       3800 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3801;
        end

       3801 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[375];
              heapArray  = localMem[409];
              ip = 3802;
              heapClock = 1;
        end

       3802 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3803;
        end

       3803 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3804;
        end

       3804 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3805;
              heapClock = 1;
        end

       3805 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3806;
        end

       3806 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1030] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3807;
              heapClock = 1;
        end

       3807 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3808;
        end

       3808 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[410] = localMem[1030];
              ip = 3809;
        end

       3809 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3810;
        end

       3810 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[375];
              heapArray  = localMem[410];
              ip = 3811;
              heapClock = 1;
        end

       3811 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3812;
        end

       3812 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[411] = localMem[400] + 1;
              ip = 3813;
        end

       3813 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1031] = localMem[411];
              ip = 3814;
        end

       3814 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3815;
        end

       3815 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[377];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1031];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3816;
              heapClock = 1;
        end

       3816 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3817;
        end

       3817 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3818;
        end

       3818 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 3819;
              heapClock = 1;
        end

       3819 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3820;
        end

       3820 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1032] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3821;
              heapClock = 1;
        end

       3821 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3822;
        end

       3822 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[412] = localMem[1032];
              ip = 3823;
        end

       3823 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1033] = localMem[378];
              ip = 3824;
        end

       3824 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3825;
        end

       3825 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[412];                                                // Array to write to
              heapIndex   = localMem[411];                                                // Index of element to write to
              heapIn      = localMem[1033];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3826;
              heapClock = 1;
        end

       3826 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3827;
        end

       3827 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4445;
        end

       3828 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3828");
        end

       3829 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3829");
        end

       3830 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  3830");
        end

       3831 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3831");
        end

       3832 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3832");
        end

       3833 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3833");
        end

       3834 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3834");
        end

       3835 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3835");
        end

       3836 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3836");
        end

       3837 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3837");
        end

       3838 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  3838");
        end

       3839 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3839");
        end

       3840 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3840");
        end

       3841 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3841");
        end

       3842 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3842");
        end

       3843 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  3843");
        end

       3844 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3844");
        end

       3845 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3845");
        end

       3846 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3846");
        end

       3847 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3847");
        end

       3848 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3848");
        end

       3849 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3849");
        end

       3850 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3850");
        end

       3851 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3851");
        end

       3852 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3852");
        end

       3853 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3853");
        end

       3854 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3854");
        end

       3855 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3855");
        end

       3856 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3856");
        end

       3857 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3857");
        end

       3858 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3858");
        end

       3859 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3859");
        end

       3860 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3860");
        end

       3861 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3861");
        end

       3862 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3862");
        end

       3863 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3863");
        end

       3864 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3864");
        end

       3865 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3865");
        end

       3866 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3866");
        end

       3867 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3867");
        end

       3868 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3868");
        end

       3869 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3869");
        end

       3870 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3870");
        end

       3871 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3871");
        end

       3872 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3872");
        end

       3873 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3873");
        end

       3874 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3874");
        end

       3875 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3875");
        end

       3876 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3876");
        end

       3877 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3877");
        end

       3878 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3878");
        end

       3879 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3879");
        end

       3880 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3880");
        end

       3881 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3881");
        end

       3882 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3882");
        end

       3883 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3883");
        end

       3884 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3884");
        end

       3885 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3885");
        end

       3886 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3886");
        end

       3887 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3887");
        end

       3888 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3888");
        end

       3889 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3889");
        end

       3890 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3890");
        end

       3891 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3891");
        end

       3892 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3892");
        end

       3893 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  3893");
        end

       3894 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3894");
        end

       3895 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3895");
        end

       3896 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3896");
        end

       3897 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3897");
        end

       3898 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3898");
        end

       3899 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3899");
        end

       3900 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3900");
        end

       3901 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3901");
        end

       3902 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  3902");
        end

       3903 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3903");
        end

       3904 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3904");
        end

       3905 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3905");
        end

       3906 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3906");
        end

       3907 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3907");
        end

       3908 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3908");
        end

       3909 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3909");
        end

       3910 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3910");
        end

       3911 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3911");
        end

       3912 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  3912");
        end

       3913 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3913");
        end

       3914 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3914");
        end

       3915 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3915");
        end

       3916 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3916");
        end

       3917 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3917");
        end

       3918 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3918");
        end

       3919 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3919");
        end

       3920 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3920");
        end

       3921 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3921");
        end

       3922 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3922");
        end

       3923 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3923");
        end

       3924 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3924");
        end

       3925 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3925");
        end

       3926 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3926");
        end

       3927 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  3927");
        end

       3928 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3928");
        end

       3929 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3929");
        end

       3930 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3930");
        end

       3931 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3931");
        end

       3932 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3932");
        end

       3933 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3933");
        end

       3934 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3934");
        end

       3935 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3935");
        end

       3936 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3936");
        end

       3937 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3937");
        end

       3938 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3938");
        end

       3939 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3939");
        end

       3940 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3940");
        end

       3941 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  3941");
        end

       3942 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3942");
        end

       3943 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3943");
        end

       3944 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3944");
        end

       3945 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3945");
        end

       3946 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3946");
        end

       3947 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3947");
        end

       3948 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3948");
        end

       3949 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3949");
        end

       3950 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3950");
        end

       3951 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  3951");
        end

       3952 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3952");
        end

       3953 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3953");
        end

       3954 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3954");
        end

       3955 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3955");
        end

       3956 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3956");
        end

       3957 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3957");
        end

       3958 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3958");
        end

       3959 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3959");
        end

       3960 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3960");
        end

       3961 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3961");
        end

       3962 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3962");
        end

       3963 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3963");
        end

       3964 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3964");
        end

       3965 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3965");
        end

       3966 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3966");
        end

       3967 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3967");
        end

       3968 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3968");
        end

       3969 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3969");
        end

       3970 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3970");
        end

       3971 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3971");
        end

       3972 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3972");
        end

       3973 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3973");
        end

       3974 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3974");
        end

       3975 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3975");
        end

       3976 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3976");
        end

       3977 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3977");
        end

       3978 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3978");
        end

       3979 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3979");
        end

       3980 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3980");
        end

       3981 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3981");
        end

       3982 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3982");
        end

       3983 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3983");
        end

       3984 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3984");
        end

       3985 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3985");
        end

       3986 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3986");
        end

       3987 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  3987");
        end

       3988 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3988");
        end

       3989 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3989");
        end

       3990 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3990");
        end

       3991 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3991");
        end

       3992 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3992");
        end

       3993 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3993");
        end

       3994 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3994");
        end

       3995 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3995");
        end

       3996 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3996");
        end

       3997 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3997");
        end

       3998 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3998");
        end

       3999 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3999");
        end

       4000 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4000");
        end

       4001 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  4001");
        end

       4002 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4002");
        end

       4003 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  4003");
        end

       4004 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4004");
        end

       4005 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4005");
        end

       4006 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4006");
        end

       4007 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4007");
        end

       4008 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4008");
        end

       4009 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4009");
        end

       4010 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4010");
        end

       4011 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  4011");
        end

       4012 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4012");
        end

       4013 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  4013");
        end

       4014 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4014");
        end

       4015 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4015");
        end

       4016 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4016");
        end

       4017 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4017");
        end

       4018 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4018");
        end

       4019 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4019");
        end

       4020 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4020");
        end

       4021 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4021");
        end

       4022 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4022");
        end

       4023 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4023");
        end

       4024 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4024");
        end

       4025 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4025");
        end

       4026 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4026");
        end

       4027 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4027");
        end

       4028 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4028");
        end

       4029 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4029");
        end

       4030 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4030");
        end

       4031 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4031");
        end

       4032 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4032");
        end

       4033 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  4033");
        end

       4034 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4034");
        end

       4035 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4035");
        end

       4036 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4036");
        end

       4037 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4037");
        end

       4038 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4038");
        end

       4039 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4039");
        end

       4040 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4040");
        end

       4041 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4041");
        end

       4042 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4042");
        end

       4043 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4043");
        end

       4044 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4044");
        end

       4045 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4045");
        end

       4046 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4046");
        end

       4047 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4047");
        end

       4048 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4048");
        end

       4049 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4049");
        end

       4050 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4050");
        end

       4051 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  4051");
        end

       4052 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  4052");
        end

       4053 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4053");
        end

       4054 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  4054");
        end

       4055 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4055");
        end

       4056 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  4056");
        end

       4057 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4057");
        end

       4058 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4058");
        end

       4059 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4059");
        end

       4060 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4060");
        end

       4061 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4061");
        end

       4062 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4062");
        end

       4063 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4063");
        end

       4064 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  4064");
        end

       4065 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4065");
        end

       4066 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  4066");
        end

       4067 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4067");
        end

       4068 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4068");
        end

       4069 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4069");
        end

       4070 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4070");
        end

       4071 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4071");
        end

       4072 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4072");
        end

       4073 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4073");
        end

       4074 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4074");
        end

       4075 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4075");
        end

       4076 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4076");
        end

       4077 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4077");
        end

       4078 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4078");
        end

       4079 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4079");
        end

       4080 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4080");
        end

       4081 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4081");
        end

       4082 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4082");
        end

       4083 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4083");
        end

       4084 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4084");
        end

       4085 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4085");
        end

       4086 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4086");
        end

       4087 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4087");
        end

       4088 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4088");
        end

       4089 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4089");
        end

       4090 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4090");
        end

       4091 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4091");
        end

       4092 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4092");
        end

       4093 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4093");
        end

       4094 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4094");
        end

       4095 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4095");
        end

       4096 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4096");
        end

       4097 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4097");
        end

       4098 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4098");
        end

       4099 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4099");
        end

       4100 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4100");
        end

       4101 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4101");
        end

       4102 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4102");
        end

       4103 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4103");
        end

       4104 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4104");
        end

       4105 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4105");
        end

       4106 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4106");
        end

       4107 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4107");
        end

       4108 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4108");
        end

       4109 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4109");
        end

       4110 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4110");
        end

       4111 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4111");
        end

       4112 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4112");
        end

       4113 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4113");
        end

       4114 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4114");
        end

       4115 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4115");
        end

       4116 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4116");
        end

       4117 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4117");
        end

       4118 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4118");
        end

       4119 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4119");
        end

       4120 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4120");
        end

       4121 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4121");
        end

       4122 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4122");
        end

       4123 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  4123");
        end

       4124 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4124");
        end

       4125 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4125");
        end

       4126 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4126");
        end

       4127 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4127");
        end

       4128 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4128");
        end

       4129 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4129");
        end

       4130 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4130");
        end

       4131 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4131");
        end

       4132 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4132");
        end

       4133 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4133");
        end

       4134 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4134");
        end

       4135 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4135");
        end

       4136 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4136");
        end

       4137 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4137");
        end

       4138 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4138");
        end

       4139 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4139");
        end

       4140 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4140");
        end

       4141 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4141");
        end

       4142 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4142");
        end

       4143 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4143");
        end

       4144 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4144");
        end

       4145 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4145");
        end

       4146 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4146");
        end

       4147 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4147");
        end

       4148 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4148");
        end

       4149 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4149");
        end

       4150 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4150");
        end

       4151 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4151");
        end

       4152 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4152");
        end

       4153 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4153");
        end

       4154 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4154");
        end

       4155 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4155");
        end

       4156 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4156");
        end

       4157 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4157");
        end

       4158 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4158");
        end

       4159 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4159");
        end

       4160 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4160");
        end

       4161 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4161");
        end

       4162 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4162");
        end

       4163 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4163");
        end

       4164 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4164");
        end

       4165 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4165");
        end

       4166 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4166");
        end

       4167 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4167");
        end

       4168 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4168");
        end

       4169 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4169");
        end

       4170 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4170");
        end

       4171 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4171");
        end

       4172 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4172");
        end

       4173 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4173");
        end

       4174 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4174");
        end

       4175 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4175");
        end

       4176 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4176");
        end

       4177 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4177");
        end

       4178 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4178");
        end

       4179 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4179");
        end

       4180 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4180");
        end

       4181 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  4181");
        end

       4182 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4182");
        end

       4183 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4183");
        end

       4184 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4184");
        end

       4185 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4185");
        end

       4186 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4186");
        end

       4187 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4187");
        end

       4188 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4188");
        end

       4189 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4189");
        end

       4190 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4190");
        end

       4191 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4191");
        end

       4192 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4192");
        end

       4193 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4193");
        end

       4194 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4194");
        end

       4195 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  4195");
        end

       4196 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4196");
        end

       4197 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4197");
        end

       4198 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4198");
        end

       4199 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4199");
        end

       4200 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4200");
        end

       4201 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4201");
        end

       4202 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4202");
        end

       4203 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4203");
        end

       4204 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4204");
        end

       4205 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  4205");
        end

       4206 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4206");
        end

       4207 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4207");
        end

       4208 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4208");
        end

       4209 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4209");
        end

       4210 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4210");
        end

       4211 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4211");
        end

       4212 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4212");
        end

       4213 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4213");
        end

       4214 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4214");
        end

       4215 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4215");
        end

       4216 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4216");
        end

       4217 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  4217");
        end

       4218 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4218");
        end

       4219 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4219");
        end

       4220 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4220");
        end

       4221 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4221");
        end

       4222 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4222");
        end

       4223 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4223");
        end

       4224 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4224");
        end

       4225 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4225");
        end

       4226 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  4226");
        end

       4227 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4227");
        end

       4228 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4228");
        end

       4229 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4229");
        end

       4230 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4230");
        end

       4231 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4231");
        end

       4232 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4232");
        end

       4233 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4233");
        end

       4234 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4234");
        end

       4235 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4235");
        end

       4236 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  4236");
        end

       4237 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4237");
        end

       4238 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4238");
        end

       4239 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4239");
        end

       4240 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4240");
        end

       4241 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4241");
        end

       4242 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4242");
        end

       4243 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4243");
        end

       4244 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4244");
        end

       4245 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4245");
        end

       4246 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4246");
        end

       4247 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4247");
        end

       4248 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  4248");
        end

       4249 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4249");
        end

       4250 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4250");
        end

       4251 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4251");
        end

       4252 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4252");
        end

       4253 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4253");
        end

       4254 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  4254");
        end

       4255 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4255");
        end

       4256 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  4256");
        end

       4257 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4257");
        end

       4258 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4258");
        end

       4259 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4259");
        end

       4260 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4260");
        end

       4261 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4261");
        end

       4262 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4262");
        end

       4263 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4263");
        end

       4264 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4264");
        end

       4265 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4265");
        end

       4266 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4266");
        end

       4267 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4267");
        end

       4268 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4268");
        end

       4269 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4269");
        end

       4270 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4270");
        end

       4271 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4271");
        end

       4272 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4272");
        end

       4273 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4273");
        end

       4274 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4274");
        end

       4275 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4275");
        end

       4276 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4276");
        end

       4277 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4277");
        end

       4278 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4278");
        end

       4279 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4279");
        end

       4280 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4280");
        end

       4281 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4281");
        end

       4282 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4282");
        end

       4283 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4283");
        end

       4284 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4284");
        end

       4285 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4285");
        end

       4286 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4286");
        end

       4287 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4287");
        end

       4288 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4288");
        end

       4289 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4289");
        end

       4290 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4290");
        end

       4291 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4291");
        end

       4292 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4292");
        end

       4293 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4293");
        end

       4294 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4294");
        end

       4295 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4295");
        end

       4296 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4296");
        end

       4297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4297");
        end

       4298 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4298");
        end

       4299 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4299");
        end

       4300 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4300");
        end

       4301 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4301");
        end

       4302 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4302");
        end

       4303 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4303");
        end

       4304 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4304");
        end

       4305 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4305");
        end

       4306 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4306");
        end

       4307 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4307");
        end

       4308 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4308");
        end

       4309 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4309");
        end

       4310 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4310");
        end

       4311 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4311");
        end

       4312 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4312");
        end

       4313 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4313");
        end

       4314 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4314");
        end

       4315 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4315");
        end

       4316 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4316");
        end

       4317 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4317");
        end

       4318 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4318");
        end

       4319 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4319");
        end

       4320 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4320");
        end

       4321 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4321");
        end

       4322 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4322");
        end

       4323 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4323");
        end

       4324 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4324");
        end

       4325 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4325");
        end

       4326 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4326");
        end

       4327 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4327");
        end

       4328 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4328");
        end

       4329 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4329");
        end

       4330 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4330");
        end

       4331 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4331");
        end

       4332 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4332");
        end

       4333 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4333");
        end

       4334 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  4334");
        end

       4335 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4335");
        end

       4336 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  4336");
        end

       4337 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4337");
        end

       4338 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4338");
        end

       4339 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4339");
        end

       4340 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4340");
        end

       4341 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4341");
        end

       4342 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4342");
        end

       4343 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4343");
        end

       4344 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4344");
        end

       4345 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4345");
        end

       4346 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4346");
        end

       4347 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4347");
        end

       4348 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4348");
        end

       4349 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4349");
        end

       4350 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4350");
        end

       4351 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4351");
        end

       4352 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4352");
        end

       4353 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4353");
        end

       4354 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4354");
        end

       4355 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4355");
        end

       4356 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4356");
        end

       4357 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4357");
        end

       4358 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4358");
        end

       4359 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4359");
        end

       4360 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4360");
        end

       4361 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4361");
        end

       4362 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4362");
        end

       4363 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4363");
        end

       4364 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4364");
        end

       4365 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4365");
        end

       4366 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4366");
        end

       4367 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4367");
        end

       4368 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4368");
        end

       4369 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4369");
        end

       4370 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4370");
        end

       4371 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4371");
        end

       4372 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4372");
        end

       4373 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4373");
        end

       4374 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4374");
        end

       4375 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4375");
        end

       4376 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4376");
        end

       4377 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4377");
        end

       4378 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4378");
        end

       4379 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4379");
        end

       4380 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4380");
        end

       4381 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4381");
        end

       4382 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4382");
        end

       4383 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4383");
        end

       4384 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4384");
        end

       4385 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4385");
        end

       4386 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4386");
        end

       4387 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4387");
        end

       4388 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4388");
        end

       4389 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4389");
        end

       4390 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4390");
        end

       4391 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4391");
        end

       4392 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4392");
        end

       4393 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4393");
        end

       4394 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4394");
        end

       4395 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4395");
        end

       4396 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4396");
        end

       4397 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4397");
        end

       4398 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4398");
        end

       4399 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4399");
        end

       4400 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4400");
        end

       4401 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4401");
        end

       4402 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4402");
        end

       4403 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4403");
        end

       4404 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4404");
        end

       4405 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4405");
        end

       4406 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4406");
        end

       4407 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4407");
        end

       4408 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4408");
        end

       4409 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4409");
        end

       4410 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4410");
        end

       4411 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4411");
        end

       4412 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4412");
        end

       4413 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4413");
        end

       4414 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4414");
        end

       4415 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4415");
        end

       4416 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4416");
        end

       4417 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4417");
        end

       4418 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4418");
        end

       4419 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4419");
        end

       4420 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4420");
        end

       4421 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4421");
        end

       4422 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4422");
        end

       4423 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  4423");
        end

       4424 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4424");
        end

       4425 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4425");
        end

       4426 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4426");
        end

       4427 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4427");
        end

       4428 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4428");
        end

       4429 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4429");
        end

       4430 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4430");
        end

       4431 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4431");
        end

       4432 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  4432");
        end

       4433 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4433");
        end

       4434 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4434");
        end

       4435 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4435");
        end

       4436 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4436");
        end

       4437 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4437");
        end

       4438 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4438");
        end

       4439 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4439");
        end

       4440 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4440");
        end

       4441 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  4441");
        end

       4442 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4442");
        end

       4443 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4443");
        end

       4444 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4444");
        end

       4445 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4446;
        end

       4446 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[371] = 1;
              ip = 4447;
        end

       4447 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4450;
        end

       4448 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4449;
        end

       4449 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[371] = 0;
              ip = 4450;
        end

       4450 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4451;
        end

       4451 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4452;
        end

       4452 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4453;
        end

       4453 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4454;
        end

       4454 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[3];
              ip = 4455;
              heapClock = 1;
        end

       4455 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4456;
        end

       4456 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1] = localMem[1] + 1;
              ip = 4457;
        end

       4457 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 27;
        end

       4458 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4459;
        end

       4459 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4460;
        end

       4460 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[478] = 0;
              ip = 4461;
        end

       4461 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4462;
        end

       4462 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[478] >= 66 ? 4647 : 4463;
        end

       4463 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4464;
        end

       4464 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 4465;
              heapClock = 1;
        end

       4465 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4466;
        end

       4466 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[479] = heapOut;
              ip = 4467;
        end

       4467 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4468;
        end

       4468 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4469;
        end

       4469 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4470;
        end

       4470 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4471;
        end

       4471 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4472;
              heapClock = 1;
        end

       4472 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4473;
        end

       4473 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1116] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4474;
              heapClock = 1;
        end

       4474 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4475;
        end

       4475 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[480] = localMem[1116];
              ip = 4476;
        end

       4476 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[480] != 0 ? 4490 : 4477;
        end

       4477 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4477");
        end

       4478 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4478");
        end

       4479 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4479");
        end

       4480 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4480");
        end

       4481 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4481");
        end

       4482 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4482");
        end

       4483 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4483");
        end

       4484 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4484");
        end

       4485 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4485");
        end

       4486 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4486");
        end

       4487 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4487");
        end

       4488 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4488");
        end

       4489 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4489");
        end

       4490 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4491;
        end

       4491 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4492;
        end

       4492 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = 0;
              ip = 4493;
        end

       4493 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4494;
        end

       4494 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[481] >= 99 ? 4614 : 4495;
        end

       4495 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4496;
        end

       4496 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4497;
              heapClock = 1;
        end

       4497 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4498;
        end

       4498 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1120] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4499;
              heapClock = 1;
        end

       4499 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4500;
        end

       4500 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[482] = localMem[1120] - 1;
              ip = 4501;
        end

       4501 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4502;
        end

       4502 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4503;
              heapClock = 1;
        end

       4503 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4504;
        end

       4504 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1121] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4505;
              heapClock = 1;
        end

       4505 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4506;
        end

       4506 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[483] = localMem[1121];
              ip = 4507;
        end

       4507 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4508;
        end

       4508 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[483];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[482];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4509;
              heapClock = 1;
        end

       4509 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4510;
        end

       4510 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1122] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4511;
              heapClock = 1;
        end

       4511 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4512;
        end

       4512 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[478] <= localMem[1122] ? 4549 : 4513;
        end

       4513 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[484] = localMem[482] + 1;
              ip = 4514;
        end

       4514 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4515;
        end

       4515 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4516;
              heapClock = 1;
        end

       4516 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4517;
        end

       4517 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1123] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4518;
              heapClock = 1;
        end

       4518 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4519;
        end

       4519 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[485] = !localMem[1123];
              ip = 4520;
        end

       4520 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[485] == 0 ? 4534 : 4521;
        end

       4521 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4521");
        end

       4522 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4522");
        end

       4523 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4523");
        end

       4524 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4524");
        end

       4525 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4525");
        end

       4526 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4526");
        end

       4527 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4527");
        end

       4528 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4528");
        end

       4529 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4529");
        end

       4530 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4530");
        end

       4531 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4531");
        end

       4532 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4532");
        end

       4533 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4533");
        end

       4534 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4535;
        end

       4535 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4536;
        end

       4536 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4537;
              heapClock = 1;
        end

       4537 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4538;
        end

       4538 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1127] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4539;
              heapClock = 1;
        end

       4539 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4540;
        end

       4540 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[486] = localMem[1127];
              ip = 4541;
        end

       4541 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4542;
        end

       4542 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[486];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[484];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4543;
              heapClock = 1;
        end

       4543 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4544;
        end

       4544 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1128] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4545;
              heapClock = 1;
        end

       4545 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4546;
        end

       4546 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[487] = localMem[1128];
              ip = 4547;
        end

       4547 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[480] = localMem[487];
              ip = 4548;
        end

       4548 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4611;
        end

       4549 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4550;
        end

       4550 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4551;
        end

       4551 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[478];
              heapAction = `Index;
              heapArray  = localMem[483];
              ip = 4552;
              heapClock = 1;
        end

       4552 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4553;
        end

       4553 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[488] = heapOut;
              ip = 4554;
        end

       4554 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4555;
        end

       4555 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4556;
        end

       4556 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[488] == 0 ? 4570 : 4557;
        end

       4557 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1129] = localMem[480];
              ip = 4558;
        end

       4558 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4559;
        end

       4559 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[479];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1129];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 4560;
              heapClock = 1;
        end

       4560 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4561;
        end

       4561 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1130] = 1;
              ip = 4562;
        end

       4562 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4563;
        end

       4563 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[479];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1130];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 4564;
              heapClock = 1;
        end

       4564 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4565;
        end

       4565 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[1131] = localMem[488] - 1;
              ip = 4566;
        end

       4566 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4567;
        end

       4567 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[479];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1131];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 4568;
              heapClock = 1;
        end

       4568 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4569;
        end

       4569 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4618;
        end

       4570 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4571;
        end

       4571 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4572;
        end

       4572 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
              heapIn     = localMem[478];
              heapAction = `Less;
              heapArray  = localMem[483];
              ip = 4573;
              heapClock = 1;
        end

       4573 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4574;
        end

       4574 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[489] = heapOut;
              ip = 4575;
        end

       4575 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4576;
        end

       4576 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4577;
        end

       4577 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4578;
        end

       4578 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4579;
              heapClock = 1;
        end

       4579 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4580;
        end

       4580 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1132] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4581;
              heapClock = 1;
        end

       4581 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4582;
        end

       4582 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[490] = !localMem[1132];
              ip = 4583;
        end

       4583 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[490] == 0 ? 4597 : 4584;
        end

       4584 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4584");
        end

       4585 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4585");
        end

       4586 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4586");
        end

       4587 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4587");
        end

       4588 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4588");
        end

       4589 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4589");
        end

       4590 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4590");
        end

       4591 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4591");
        end

       4592 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4592");
        end

       4593 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4593");
        end

       4594 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4594");
        end

       4595 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4595");
        end

       4596 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4596");
        end

       4597 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4598;
        end

       4598 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4599;
        end

       4599 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4600;
              heapClock = 1;
        end

       4600 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4601;
        end

       4601 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1136] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4602;
              heapClock = 1;
        end

       4602 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4603;
        end

       4603 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[491] = localMem[1136];
              ip = 4604;
        end

       4604 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4605;
        end

       4605 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[491];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[489];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4606;
              heapClock = 1;
        end

       4606 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4607;
        end

       4607 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1137] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4608;
              heapClock = 1;
        end

       4608 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4609;
        end

       4609 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[492] = localMem[1137];
              ip = 4610;
        end

       4610 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[480] = localMem[492];
              ip = 4611;
        end

       4611 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4612;
        end

       4612 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[481] = localMem[481] + 1;
              ip = 4613;
        end

       4613 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4493;
        end

       4614 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4614");
        end

       4615 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  4615");
        end

       4616 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4616");
        end

       4617 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4617");
        end

       4618 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4619;
        end

       4619 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4620;
        end

       4620 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[479];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4621;
              heapClock = 1;
        end

       4621 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4622;
        end

       4622 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1138] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4623;
              heapClock = 1;
        end

       4623 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4624;
        end

       4624 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[493] = localMem[1138];
              ip = 4625;
        end

       4625 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4626;
        end

       4626 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[479];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4627;
              heapClock = 1;
        end

       4627 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4628;
        end

       4628 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1139] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4629;
              heapClock = 1;
        end

       4629 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4630;
        end

       4630 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[494] = localMem[1139];
              ip = 4631;
        end

       4631 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4632;
        end

       4632 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[493];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4633;
              heapClock = 1;
        end

       4633 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4634;
        end

       4634 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1140] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4635;
              heapClock = 1;
        end

       4635 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4636;
        end

       4636 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[495] = localMem[1140];
              ip = 4637;
        end

       4637 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4638;
        end

       4638 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[495];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[494];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4639;
              heapClock = 1;
        end

       4639 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4640;
        end

       4640 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1141] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4641;
              heapClock = 1;
        end

       4641 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4642;
        end

       4642 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[496] = localMem[1141];
              ip = 4643;
        end

       4643 :
        begin                                                                   // out
          //$display("AAAA %4d %4d out", steps, ip);
              outMem[outMemPos] = localMem[496];
              outMemPos = outMemPos + 1;
              ip = 4644;
        end

       4644 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4645;
        end

       4645 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[478] = localMem[478] + 1;
              ip = 4646;
        end

       4646 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4461;
        end

       4647 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4648;
        end

       4648 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4649;
        end

       4649 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 4650;
              heapClock = 1;
        end

       4650 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4651;
        end

       4651 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[497] = heapOut;
              ip = 4652;
        end

       4652 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4653;
        end

       4653 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4654;
        end

       4654 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4655;
        end

       4655 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4656;
        end

       4656 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4657;
              heapClock = 1;
        end

       4657 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4658;
        end

       4658 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1142] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4659;
              heapClock = 1;
        end

       4659 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4660;
        end

       4660 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[498] = localMem[1142];
              ip = 4661;
        end

       4661 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[498] != 0 ? 4675 : 4662;
        end

       4662 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4662");
        end

       4663 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4663");
        end

       4664 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4664");
        end

       4665 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4665");
        end

       4666 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4666");
        end

       4667 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4667");
        end

       4668 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4668");
        end

       4669 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4669");
        end

       4670 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4670");
        end

       4671 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4671");
        end

       4672 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4672");
        end

       4673 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4673");
        end

       4674 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4674");
        end

       4675 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4676;
        end

       4676 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4677;
        end

       4677 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[499] = 0;
              ip = 4678;
        end

       4678 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4679;
        end

       4679 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[499] >= 99 ? 4799 : 4680;
        end

       4680 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4681;
        end

       4681 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4682;
              heapClock = 1;
        end

       4682 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4683;
        end

       4683 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1146] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4684;
              heapClock = 1;
        end

       4684 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4685;
        end

       4685 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[500] = localMem[1146] - 1;
              ip = 4686;
        end

       4686 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4687;
        end

       4687 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4688;
              heapClock = 1;
        end

       4688 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4689;
        end

       4689 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1147] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4690;
              heapClock = 1;
        end

       4690 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4691;
        end

       4691 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[501] = localMem[1147];
              ip = 4692;
        end

       4692 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4693;
        end

       4693 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[501];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[500];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4694;
              heapClock = 1;
        end

       4694 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4695;
        end

       4695 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1148] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4696;
              heapClock = 1;
        end

       4696 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4697;
        end

       4697 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = 66 <= localMem[1148] ? 4734 : 4698;
        end

       4698 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[502] = localMem[500] + 1;
              ip = 4699;
        end

       4699 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4700;
        end

       4700 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4701;
              heapClock = 1;
        end

       4701 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4702;
        end

       4702 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1149] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4703;
              heapClock = 1;
        end

       4703 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4704;
        end

       4704 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[503] = !localMem[1149];
              ip = 4705;
        end

       4705 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[503] == 0 ? 4719 : 4706;
        end

       4706 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1150] = localMem[498];
              ip = 4707;
        end

       4707 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4708;
        end

       4708 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[497];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1150];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 4709;
              heapClock = 1;
        end

       4709 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4710;
        end

       4710 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1151] = 2;
              ip = 4711;
        end

       4711 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4712;
        end

       4712 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[497];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1151];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 4713;
              heapClock = 1;
        end

       4713 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4714;
        end

       4714 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1152] = localMem[502];
              ip = 4715;
        end

       4715 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4716;
        end

       4716 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[497];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1152];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 4717;
              heapClock = 1;
        end

       4717 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4718;
        end

       4718 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4803;
        end

       4719 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4720;
        end

       4720 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4721;
        end

       4721 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4722;
              heapClock = 1;
        end

       4722 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4723;
        end

       4723 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1153] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4724;
              heapClock = 1;
        end

       4724 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4725;
        end

       4725 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[504] = localMem[1153];
              ip = 4726;
        end

       4726 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4727;
        end

       4727 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[504];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[502];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4728;
              heapClock = 1;
        end

       4728 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4729;
        end

       4729 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1154] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4730;
              heapClock = 1;
        end

       4730 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4731;
        end

       4731 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[505] = localMem[1154];
              ip = 4732;
        end

       4732 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[498] = localMem[505];
              ip = 4733;
        end

       4733 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4796;
        end

       4734 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4734");
        end

       4735 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4735");
        end

       4736 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  4736");
        end

       4737 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4737");
        end

       4738 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  4738");
        end

       4739 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4739");
        end

       4740 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4740");
        end

       4741 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  4741");
        end

       4742 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4742");
        end

       4743 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4743");
        end

       4744 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4744");
        end

       4745 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4745");
        end

       4746 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4746");
        end

       4747 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4747");
        end

       4748 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4748");
        end

       4749 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4749");
        end

       4750 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  4750");
        end

       4751 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4751");
        end

       4752 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4752");
        end

       4753 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4753");
        end

       4754 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4754");
        end

       4755 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4755");
        end

       4756 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4756");
        end

       4757 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed  4757");
        end

       4758 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4758");
        end

       4759 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  4759");
        end

       4760 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4760");
        end

       4761 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4761");
        end

       4762 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4762");
        end

       4763 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4763");
        end

       4764 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4764");
        end

       4765 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4765");
        end

       4766 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4766");
        end

       4767 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  4767");
        end

       4768 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  4768");
        end

       4769 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4769");
        end

       4770 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4770");
        end

       4771 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4771");
        end

       4772 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4772");
        end

       4773 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4773");
        end

       4774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4774");
        end

       4775 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4775");
        end

       4776 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4776");
        end

       4777 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4777");
        end

       4778 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4778");
        end

       4779 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  4779");
        end

       4780 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4780");
        end

       4781 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  4781");
        end

       4782 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4782");
        end

       4783 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4783");
        end

       4784 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4784");
        end

       4785 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4785");
        end

       4786 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4786");
        end

       4787 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4787");
        end

       4788 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4788");
        end

       4789 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4789");
        end

       4790 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  4790");
        end

       4791 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4791");
        end

       4792 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  4792");
        end

       4793 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  4793");
        end

       4794 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4794");
        end

       4795 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  4795");
        end

       4796 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4797;
        end

       4797 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[499] = localMem[499] + 1;
              ip = 4798;
        end

       4798 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 4678;
        end

       4799 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4799");
        end

       4800 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  4800");
        end

       4801 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4801");
        end

       4802 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  4802");
        end

       4803 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 4804;
        end

       4804 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4805;
        end

       4805 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[497];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                               // Request a read, not a write
              ip = 4806;
              heapClock = 1;
        end

       4806 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4807;
        end

       4807 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1164] = heapOut;                                                     // Data retrieved from heap memory
              ip = 4808;
              heapClock = 1;
        end

       4808 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 4809;
        end

       4809 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[511] = localMem[1164];
              ip = 4810;
        end

       4810 :
        begin                                                                   // out
          //$display("AAAA %4d %4d out", steps, ip);
              outMem[outMemPos] = localMem[511];
              outMemPos = outMemPos + 1;
              ip = 4811;
        end
      endcase
      success = outMem[0] == 0 && outMem[1] == 2 && outMem[2] == 4 && outMem[3] == 6 && outMem[4] == 8 && outMem[5] == 10 && outMem[6] == 12 && outMem[7] == 14 && outMem[8] == 16 && outMem[9] == 18 && outMem[10] == 20 && outMem[11] == 22 && outMem[12] == 24 && outMem[13] == 26 && outMem[14] == 28 && outMem[15] == 30 && outMem[16] == 32 && outMem[17] == 34 && outMem[18] == 36 && outMem[19] == 38 && outMem[20] == 40 && outMem[21] == 42 && outMem[22] == 44 && outMem[23] == 46 && outMem[24] == 48 && outMem[25] == 50 && outMem[26] == 52 && outMem[27] == 54 && outMem[28] == 56 && outMem[29] == 58 && outMem[30] == 60 && outMem[31] == 62 && outMem[32] == 64 && outMem[33] == 66 && outMem[34] == 68 && outMem[35] == 70 && outMem[36] == 72 && outMem[37] == 74 && outMem[38] == 76 && outMem[39] == 78 && outMem[40] == 80 && outMem[41] == 82 && outMem[42] == 84 && outMem[43] == 86 && outMem[44] == 88 && outMem[45] == 90 && outMem[46] == 92 && outMem[47] == 94 && outMem[48] == 96 && outMem[49] == 98 && outMem[50] == 100 && outMem[51] == 102 && outMem[52] == 104 && outMem[53] == 106 && outMem[54] == 108 && outMem[55] == 110 && outMem[56] == 112 && outMem[57] == 114 && outMem[58] == 116 && outMem[59] == 118 && outMem[60] == 120 && outMem[61] == 122 && outMem[62] == 124 && outMem[63] == 126 && outMem[64] == 128 && outMem[65] == 130 && outMem[66] == 2;
      steps = steps + 1;
      finished = steps >  62704;
    end
  end

endmodule
