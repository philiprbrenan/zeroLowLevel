// Check double frees, over allocation
// Check access to unallocated arrays or elements
// Check push overflow, pop underflow
// Next Message 10000280
`define Reset        1  /* Zero all memory sizes                               */
`define Write        2  /* Write an element                                    */
`define Read         3  /* Read an element                                     */
`define Size         4  /* Size of array                                       */
`define Inc          5  /* Increment size of array if possible                 */
`define Dec          6  /* Decrement size of array if possible                 */
`define Index        7  /* Index of element in array                           */
`define Less         8  /* Elements of array less than in                      */
`define Greater      9  /* Elements of array greater than in                   */
`define Up          10  /* Move array up                                       */
`define Down        11  /* Move array down                                     */
`define Long1       12  /* Move long first step                                */
`define Long2       13  /* Move long last  step                                */
`define Push        14  /* Push if possible                                    */
`define Pop         15  /* Pop if possible                                     */
`define Dump        16  /* Dump                                                */
`define Resize      17  /* Resize an array                                     */
`define Alloc       18  /* Allocate a new array before using it                */
`define Free        19  /* Free an array for reuse                             */
`define Add         20  /* Add to an element returning the new value           */
`define AddAfter    21  /* Add to an element returning the previous value      */
`define Subtract    22  /* Subtract to an element returning the new value      */
`define SubAfter    23  /* Subtract to an element returning the previous value */
`define ShiftLeft   24  /* Shift left                                          */
`define ShiftRight  25  /* Shift right                                         */
`define NotLogical  26  /* Not - logical                                       */
`define Not         27  /* Not - bitwise                                       */
`define Or          28  /* Or                                                  */
`define Xor         29  /* Xor                                                 */
`define And         30  /* And                                                 */

module Memory
#(parameter integer ADDRESS_BITS =  8,                                          // Number of bits in an address
  parameter integer INDEX_BITS   =  3,                                          // Bits in in an index
  parameter integer DATA_BITS    = 16)                                          // Width of an element in bits
 (input wire                    clock,                                          // Clock to drive array operations
  input wire[7:0]               action,                                         // Operation to be performed on array
  input wire [ADDRESS_BITS-1:0] array,                                          // The number of the array to work on
  input wire [INDEX_BITS  -1:0] index,                                          // Index within array
  input wire [DATA_BITS   -1:0] in,                                             // Input data
  output reg [DATA_BITS   -1:0] out,                                            // Output data
  output reg [31:0]             error);                                         // Error

  parameter integer ARRAY_LENGTH = 2**INDEX_BITS;                               // Maximum index
  parameter integer ARRAYS       = 2**ADDRESS_BITS;                             // Number of memory elements for both arrays and elements

  reg [DATA_BITS   -1:0] memory     [ARRAYS-1:0][ARRAY_LENGTH-1:0];             // Memory containing arrays in fixed blocks
  reg [DATA_BITS   -1:0] copy                   [ARRAY_LENGTH-1:0];             // Copy of one array
  reg [INDEX_BITS    :0] arraySizes [ARRAYS-1:0];                               // Current size of each array
  reg [ADDRESS_BITS-1:0] freedArrays[ARRAYS-1:0];                               // Currently freed arrays
  reg                    allocations[ARRAYS-1:0];                               // Currently allocated arrays

  integer allocatedArrays;                                                      // Arrays allocated
  integer freedArraysTop;                                                       // Top of the freed arrays stack
  integer result;                                                               // Result of each array operation
  integer size;                                                                 // Size of current array
  integer moveLongStartArray;                                                   // Source array of move long
  integer moveLongStartIndex;                                                   // Source index of move long
  integer i, a, b;                                                              // Index

  task checkWriteable(input integer err);                                       // Check a memory is writable
    begin
       error = 0;
       if (array >= allocatedArrays) begin
         //$display("Array has not been allocated, array %d", array);
         error = err;
       end
       if (!allocations[array]) begin
         //$display("Array has been freed, array %d", array);
         error = err + 1;
       end
    end
  endtask

  task checkReadable(input integer err);                                        // Check a memory locationis readable
    begin
       checkWriteable(err);
       if (index >= arraySizes[array]) begin
         //$display("Access outside array bounds, array %d, size: %d, access: %d", array, arraySizes[array], index);
         error = err + 2;
       end
    end
  endtask

  task dump;                                                                    // Dump some memory
    begin
      //$display("    %2d %2d %2d", arraySizes[0], arraySizes[1], arraySizes[2]);
      for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
        //$display("%2d  %2d %2d %2d", i, memory[0][i], memory[1][i], memory[2][i]);
      end
    end
  endtask

  always @(clock) begin                                                             // Each transition
    case(action)                                                                // Decode request
      `Reset: begin                                                             // Reset
        freedArraysTop = 0;                                                     // Free all arrays
        allocatedArrays = 0;
      end

      `Write: begin                                                             // Write
        checkWriteable(10000010);
        if (!error) begin
          memory[array][index] = in;
          if (index >= arraySizes[array] && index < ARRAY_LENGTH) begin
            arraySizes[array] = index + 1;
          end
          out = in;
        end
      end

      `Read: begin                                                              // Read
        checkReadable(10000020);
        if (!error) begin
          out = memory[array][index];
        end
      end

      `Size: begin                                                              // Size
        checkWriteable(10000030);
        if (!error) begin
          out = arraySizes[array];
        end
      end

      `Dec: begin                                                               // Decrement
        checkWriteable(10000040);
        if (!error) begin
          if (arraySizes[array] > 0) arraySizes[array] = arraySizes[array] - 1;
          else begin
            //$display("Attempt to decrement empty array, array %d", array); error = 10000044;
          end
        end
      end

      `Inc: begin                                                               // Increment
        checkWriteable(10000050);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;
          else begin
            //$display("Attempt to decrement full array, array %d", array);  error = 10000054;
          end
        end
      end

      `Index: begin                                                             // Index
        checkWriteable(10000060);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] == in) result = i + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Less: begin                                                              // Count less
        checkWriteable(10000070);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] < in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Greater: begin                                                           // Count greater
        checkWriteable(10000080);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] > in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Down: begin                                                              // Down
        checkWriteable(10000270);
        if (!error) begin
          size   = arraySizes[array];
          if (size > 0) begin
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i]; // Copy source array
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                       // Move original array up
              if (i > index && i <= size) begin
                memory[array][i-1] = copy[i];
              end
            end
            out = copy[index];                                                  // Return replaced value
            arraySizes[array] = arraySizes[array] - 1;                          // Decrease array size
          end
          else error = 100000274;                                               // Orignal array was emoty so we cannot shift it down
        end
      end

      `Up: begin                                                                // Up
        checkWriteable(10000090);
        if (!error) begin
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i];   // Copy source array
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Move original array up
            if (i > index && i <= size) begin
              memory[array][i] = copy[i-1];
            end
          end
          memory[array][index] = in;                                            // Insert new value
          if (size < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;   // Increase array size
        end
      end

      `Long1: begin                                                             // Move long start
        checkReadable(10000100);
        if (!error) begin
          moveLongStartArray = array;                                           // Record source
          moveLongStartIndex = index;
        end
      end

      `Long2: begin                                                             // Move long finish
        checkWriteable(10000110);
        if (!error) begin
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Copy from source to target
            if (i < in && index + i < ARRAY_LENGTH && moveLongStartIndex+i < ARRAY_LENGTH) begin
              memory[array][index+i] = memory[moveLongStartArray][moveLongStartIndex+i];
              if (index+i >= arraySizes[array]) arraySizes[array] = index+i+1;
            end
          end
        end
      end

      `Push: begin                                                              // Push
        checkWriteable(10000120);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) begin
            memory[array][arraySizes[array]] = in;
            arraySizes[array] = arraySizes[array] + 1;
          end
          else begin
            //$display("Attempt to push to full array, array %d, value %d", array, in);  error = 10000124;
          end
        end
      end

      `Pop: begin                                                               // Pop
        checkWriteable(10000130);
        if (!error) begin
          if (arraySizes[array] > 0) begin
            arraySizes[array] = arraySizes[array] - 1;
            out = memory[array][arraySizes[array]];
          end
          else begin
            //$display("Attempt to pop empty array, array %d", array); error = 10000134;
          end
        end
      end

      `Dump: begin                                                              // Dump
        dump();
      end

      `Resize: begin                                                            // Resize
        checkWriteable(10000140);
        if (!error) begin
          if (in <= ARRAY_LENGTH) arraySizes[array] = in;
          else begin
            //$display("Attempt to make an array too large, array %d, max %d, size %d", array, ARRAY_LENGTH, in); error = 10000144;
          end
        end
      end

      `Alloc: begin                                                             // Allocate an array
        if (freedArraysTop > 0) begin                                           // Reuse a freed array
          freedArraysTop = freedArraysTop - 1;
          result = freedArrays[freedArraysTop];
        end
        else if (allocatedArrays < ARRAYS-1) begin                              // Allocate a new array - assumes enough memory
          result          = allocatedArrays;
          allocatedArrays = allocatedArrays + 1;
        end
        else begin
          //$display("Out of memory, cannot allocate a new array"); error = 10000270;
        end
        allocations[result] = 1;                                                // Allocated
        arraySizes[result] = 0;                                                 // Empty array
        out = result;
      end

      `Free: begin                                                              // Free an array
        checkWriteable(10000150);
        if (!error) begin
          freedArrays[freedArraysTop] = array;                                  // Relies on the user not re freeing a freed array - we should probably hve another array to prevent this
          allocations[freedArraysTop] = 0;                                      // No longer allocated
          freedArraysTop = freedArraysTop + 1;
        end
      end

      `Add: begin                                                               // Add to an element
        checkReadable(10000160);
        if (!error) begin
          memory[array][index] = memory[array][index] + in;
          out = memory[array][index];
        end
      end

      `AddAfter: begin                                                          // Add to an element after putting the content of the element on out
        checkReadable(10000170);
        if (!error) begin
        out = memory[array][index];
        memory[array][index] = memory[array][index] + in;
        end
      end

      `Subtract: begin                                                          // Subtract from an element
        checkReadable(10000180);
        if (!error) begin
          memory[array][index] = memory[array][index] - in;
          out = memory[array][index];
        end
      end

      `SubAfter: begin                                                          // Subtract from an element after putting the content of the element on out
        checkReadable(10000190);
        if (!error) begin
          out = memory[array][index];
          memory[array][index] = memory[array][index] - in;
        end
      end

      `ShiftLeft: begin                                                         // Shift left
        checkReadable(10000200);
        if (!error) begin
          memory[array][index] = memory[array][index] << in;
          out = memory[array][index];
        end
      end

      `ShiftRight: begin                                                        // Shift right
        checkReadable(10000210);
        if (!error) begin
          memory[array][index] = memory[array][index] >> in;
          out = memory[array][index];
        end
      end

      `NotLogical: begin                                                        // Not logical
        checkReadable(10000220);
        if (!error) begin
          memory[array][index] = !memory[array][index];
          out = memory[array][index];
        end
      end

      `Not: begin                                                               // Not
        checkReadable(10000230);
        if (!error) begin
          memory[array][index] = ~memory[array][index];
          out = memory[array][index];
        end
      end

      `Or: begin                                                                // Or
        checkReadable(10000240);
        if (!error) begin
          memory[array][index] = memory[array][index] | in;
          out = memory[array][index];
        end
      end

      `Xor: begin                                                               // Xor
        checkReadable(10000250);
        if (!error) begin
          memory[array][index] = memory[array][index] ^ in;
          out = memory[array][index];
        end
      end

      `And: begin                                                               // And
        checkReadable(10000260);
        if (!error) begin
          memory[array][index] = memory[array][index] & in;
          out = memory[array][index];
        end
      end
    endcase
  end
endmodule
//-----------------------------------------------------------------------------
// Fpga test
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga                                                                     // Run test programs
 (input  wire clock,                                                            // Driving clock
  input  wire reset,                                                            // Restart program
  output reg  finished,                                                         // Goes high when the program has finished
  output reg  success);                                                         // Goes high on finish if all the tests passed

  reg                heapClock;                                                 // Clock to drive array operations
  reg [7:0]          heapAction;                                                // Operation to be performed on array
  reg [       9-1:0] heapArray;                                         // The number of the array to work on
  reg [       3-1:0] heapIndex;                                         // Index within array
  reg [      12-1:0] heapIn;                                            // Input data
  reg [      12-1:0] heapOut;                                           // Output data
  reg [31        :0] heapError;                                                 // Error on heap operation if not zero

  Memory                                                                        // Memory module
   #(       9,        3,       12)                          // Address bits, index bits, data bits
    heap(                                                                       // Create heap memory
    .clock  (heapClock),
    .action (heapAction),
    .array  (heapArray),
    .index  (heapIndex),
    .in     (heapIn),
    .out    (heapOut),
    .error  (heapError)
  );
  reg [      12-1:0] localMem[    1204-1:0];                       // Local memory
  reg [      12-1:0]   outMem[       1  -1:0];                       // Out channel
  reg [      12-1:0]    inMem[       1   -1:0];                       // In channel

  integer inMemPos;                                                             // Current position in input channel
  integer outMemPos;                                                            // Position in output channel

  integer ip;                                                                   // Instruction pointer
  integer steps;                                                                // Number of steps executed so far
  integer i, j, k;                                                              // A useful counter

  always @(posedge clock, negedge clock) begin                                  // Each instruction
    if (reset) begin
      ip             = 0;
      steps          = 0;
      inMemPos       = 0;
      outMemPos      = 0;
      finished       = 0;
      success        = 0;

    end
    else begin
      steps = steps + 1;
      case(ip)

          0 :
        begin                                                                   // start
          //$display("AAAA %4d %4d start", steps, ip);
              heapClock = 0;                                                    // Ready for next operation
              ip = 1;
        end

          1 :
        begin                                                                   // start2
          //$display("AAAA %4d %4d start2", steps, ip);
              heapAction = `Reset;                                          // Ready for next operation
              ip = 2;
              heapClock = ~ heapClock;
        end

          2 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3;
              heapClock = ~ heapClock;
        end

          3 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[0] = heapOut;
              ip = 4;
        end

          4 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[528] = 3;
              ip = 5;
        end

          5 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[528];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 6;
              heapClock = ~ heapClock;
        end

          6 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[529] = 0;
              ip = 7;
        end

          7 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[529];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 8;
              heapClock = ~ heapClock;
        end

          8 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[530] = 0;
              ip = 9;
        end

          9 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[530];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 10;
              heapClock = ~ heapClock;
        end

         10 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[531] = 0;
              ip = 11;
        end

         11 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[531];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 12;
              heapClock = ~ heapClock;
        end

         12 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 13;
        end

         13 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1] = 0;
              ip = 14;
        end

         14 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 15;
        end

         15 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[1] >= 66 ? 2189 : 16;
        end

         16 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[2] = localMem[1] + localMem[1];
              ip = 17;
        end

         17 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 18;
              heapClock = ~ heapClock;
        end

         18 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[3] = heapOut;
              ip = 19;
        end

         19 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 20;
        end

         20 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 21;
              heapClock = ~ heapClock;
        end

         21 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[532] = heapOut;                                                     // Data retrieved from heap memory
              ip = 22;
              heapClock = ~ heapClock;
        end

         22 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[4] = localMem[532];
              ip = 23;
        end

         23 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[4] != 0 ? 75 : 24;
        end

         24 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 25;
              heapClock = ~ heapClock;
        end

         25 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[5] = heapOut;
              ip = 26;
        end

         26 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[533] = 1;
              ip = 27;
        end

         27 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[533];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 28;
              heapClock = ~ heapClock;
        end

         28 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[534] = 0;
              ip = 29;
        end

         29 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[534];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 30;
              heapClock = ~ heapClock;
        end

         30 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 31;
              heapClock = ~ heapClock;
        end

         31 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[6] = heapOut;
              ip = 32;
        end

         32 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[535] = localMem[6];
              ip = 33;
        end

         33 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[535];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 34;
              heapClock = ~ heapClock;
        end

         34 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 35;
              heapClock = ~ heapClock;
        end

         35 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[7] = heapOut;
              ip = 36;
        end

         36 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[536] = localMem[7];
              ip = 37;
        end

         37 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[536];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 38;
              heapClock = ~ heapClock;
        end

         38 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[537] = 0;
              ip = 39;
        end

         39 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[537];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 40;
              heapClock = ~ heapClock;
        end

         40 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[538] = localMem[0];
              ip = 41;
        end

         41 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[538];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 42;
              heapClock = ~ heapClock;
        end

         42 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 43;
              heapClock = ~ heapClock;
        end

         43 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[539] = heapOut;                                                     // Data retrieved from heap memory
              ip = 44;
              heapClock = ~ heapClock;
        end

         44 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[540] = localMem[539] + 1;
              ip = 45;
        end

         45 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[540];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 46;
              heapClock = ~ heapClock;
        end

         46 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 47;
              heapClock = ~ heapClock;
        end

         47 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[541] = heapOut;                                                     // Data retrieved from heap memory
              ip = 48;
              heapClock = ~ heapClock;
        end

         48 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[542] = localMem[541];
              ip = 49;
        end

         49 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[542];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 50;
              heapClock = ~ heapClock;
        end

         50 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 51;
              heapClock = ~ heapClock;
        end

         51 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[543] = heapOut;                                                     // Data retrieved from heap memory
              ip = 52;
              heapClock = ~ heapClock;
        end

         52 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[8] = localMem[543];
              ip = 53;
        end

         53 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[544] = localMem[1];
              ip = 54;
        end

         54 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[8];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[544];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 55;
              heapClock = ~ heapClock;
        end

         55 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 56;
              heapClock = ~ heapClock;
        end

         56 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[545] = heapOut;                                                     // Data retrieved from heap memory
              ip = 57;
              heapClock = ~ heapClock;
        end

         57 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[9] = localMem[545];
              ip = 58;
        end

         58 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[546] = localMem[2];
              ip = 59;
        end

         59 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[9];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[546];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 60;
              heapClock = ~ heapClock;
        end

         60 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 61;
              heapClock = ~ heapClock;
        end

         61 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[547] = heapOut;                                                     // Data retrieved from heap memory
              ip = 62;
              heapClock = ~ heapClock;
        end

         62 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[548] = localMem[547] + 1;
              ip = 63;
        end

         63 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[548];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 64;
              heapClock = ~ heapClock;
        end

         64 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[549] = localMem[5];
              ip = 65;
        end

         65 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[549];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 66;
              heapClock = ~ heapClock;
        end

         66 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 67;
              heapClock = ~ heapClock;
        end

         67 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[550] = heapOut;                                                     // Data retrieved from heap memory
              ip = 68;
              heapClock = ~ heapClock;
        end

         68 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[10] = localMem[550];
              ip = 69;
        end

         69 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[10];
              ip = 70;
              heapClock = ~ heapClock;
        end

         70 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 71;
              heapClock = ~ heapClock;
        end

         71 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[551] = heapOut;                                                     // Data retrieved from heap memory
              ip = 72;
              heapClock = ~ heapClock;
        end

         72 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[11] = localMem[551];
              ip = 73;
        end

         73 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[11];
              ip = 74;
              heapClock = ~ heapClock;
        end

         74 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2184;
        end

         75 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 76;
        end

         76 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 77;
              heapClock = ~ heapClock;
        end

         77 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[552] = heapOut;                                                     // Data retrieved from heap memory
              ip = 78;
              heapClock = ~ heapClock;
        end

         78 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[12] = localMem[552];
              ip = 79;
        end

         79 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 80;
              heapClock = ~ heapClock;
        end

         80 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[553] = heapOut;                                                     // Data retrieved from heap memory
              ip = 81;
              heapClock = ~ heapClock;
        end

         81 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[13] = localMem[553];
              ip = 82;
        end

         82 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[12] >= localMem[13] ? 152 : 83;
        end

         83 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 84;
              heapClock = ~ heapClock;
        end

         84 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[554] = heapOut;                                                     // Data retrieved from heap memory
              ip = 85;
              heapClock = ~ heapClock;
        end

         85 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[14] = localMem[554];
              ip = 86;
        end

         86 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[14] != 0 ? 151 : 87;
        end

         87 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 88;
              heapClock = ~ heapClock;
        end

         88 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[555] = heapOut;                                                     // Data retrieved from heap memory
              ip = 89;
              heapClock = ~ heapClock;
        end

         89 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[15] = !localMem[555];
              ip = 90;
        end

         90 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[15] == 0 ? 150 : 91;
        end

         91 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 92;
              heapClock = ~ heapClock;
        end

         92 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[556] = heapOut;                                                     // Data retrieved from heap memory
              ip = 93;
              heapClock = ~ heapClock;
        end

         93 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[16] = localMem[556];
              ip = 94;
        end

         94 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[1];
              heapAction = `Index;
              heapArray  = localMem[16];
              ip = 95;
              heapClock = ~ heapClock;
        end

         95 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[17] = heapOut;
              ip = 96;
        end

         96 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[17] == 0 ? 104 : 97;
        end

         97 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed    97");
        end

         98 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed    98");
        end

         99 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed    99");
        end

        100 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   100");
        end

        101 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   101");
        end

        102 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   102");
        end

        103 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   103");
        end

        104 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 105;
        end

        105 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[12];
              heapArray  = localMem[16];
              ip = 106;
              heapClock = ~ heapClock;
        end

        106 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 107;
              heapClock = ~ heapClock;
        end

        107 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[559] = heapOut;                                                     // Data retrieved from heap memory
              ip = 108;
              heapClock = ~ heapClock;
        end

        108 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[19] = localMem[559];
              ip = 109;
        end

        109 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[12];
              heapArray  = localMem[19];
              ip = 110;
              heapClock = ~ heapClock;
        end

        110 :
        begin                                                                   // arrayCountGreater
          //$display("AAAA %4d %4d arrayCountGreater", steps, ip);
              heapIn     = localMem[1];
              heapAction = `Greater;
              heapArray  = localMem[16];
              ip = 111;
              heapClock = ~ heapClock;
        end

        111 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[20] = heapOut;
              ip = 112;
        end

        112 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[20] != 0 ? 130 : 113;
        end

        113 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 114;
              heapClock = ~ heapClock;
        end

        114 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[560] = heapOut;                                                     // Data retrieved from heap memory
              ip = 115;
              heapClock = ~ heapClock;
        end

        115 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[21] = localMem[560];
              ip = 116;
        end

        116 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[561] = localMem[1];
              ip = 117;
        end

        117 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[21];                                                // Array to write to
              heapIndex   = localMem[12];                                                // Index of element to write to
              heapIn      = localMem[561];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 118;
              heapClock = ~ heapClock;
        end

        118 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 119;
              heapClock = ~ heapClock;
        end

        119 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[562] = heapOut;                                                     // Data retrieved from heap memory
              ip = 120;
              heapClock = ~ heapClock;
        end

        120 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[22] = localMem[562];
              ip = 121;
        end

        121 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[563] = localMem[2];
              ip = 122;
        end

        122 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[22];                                                // Array to write to
              heapIndex   = localMem[12];                                                // Index of element to write to
              heapIn      = localMem[563];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 123;
              heapClock = ~ heapClock;
        end

        123 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[564] = localMem[12] + 1;
              ip = 124;
        end

        124 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[4];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[564];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 125;
              heapClock = ~ heapClock;
        end

        125 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 126;
              heapClock = ~ heapClock;
        end

        126 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[565] = heapOut;                                                     // Data retrieved from heap memory
              ip = 127;
              heapClock = ~ heapClock;
        end

        127 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[566] = localMem[565] + 1;
              ip = 128;
        end

        128 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[566];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 129;
              heapClock = ~ heapClock;
        end

        129 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2184;
        end

        130 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   130");
        end

        131 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed   131");
        end

        132 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   132");
        end

        133 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   133");
        end

        134 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   134");
        end

        135 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   135");
        end

        136 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   136");
        end

        137 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   137");
        end

        138 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   138");
        end

        139 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   139");
        end

        140 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   140");
        end

        141 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   141");
        end

        142 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   142");
        end

        143 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   143");
        end

        144 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   144");
        end

        145 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   145");
        end

        146 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   146");
        end

        147 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   147");
        end

        148 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   148");
        end

        149 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   149");
        end

        150 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 151;
        end

        151 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 152;
        end

        152 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 153;
        end

        153 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 154;
              heapClock = ~ heapClock;
        end

        154 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[573] = heapOut;                                                     // Data retrieved from heap memory
              ip = 155;
              heapClock = ~ heapClock;
        end

        155 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[26] = localMem[573];
              ip = 156;
        end

        156 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 157;
        end

        157 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 158;
              heapClock = ~ heapClock;
        end

        158 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[574] = heapOut;                                                     // Data retrieved from heap memory
              ip = 159;
              heapClock = ~ heapClock;
        end

        159 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[28] = localMem[574];
              ip = 160;
        end

        160 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 161;
              heapClock = ~ heapClock;
        end

        161 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[575] = heapOut;                                                     // Data retrieved from heap memory
              ip = 162;
              heapClock = ~ heapClock;
        end

        162 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[29] = localMem[575];
              ip = 163;
        end

        163 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 164;
              heapClock = ~ heapClock;
        end

        164 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[576] = heapOut;                                                     // Data retrieved from heap memory
              ip = 165;
              heapClock = ~ heapClock;
        end

        165 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[30] = localMem[576];
              ip = 166;
        end

        166 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[28] <  localMem[30] ? 626 : 167;
        end

        167 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[31] = localMem[30];
              ip = 168;
        end

        168 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[31] = localMem[31] >> 1;
              ip = 169;
              ip = 169;
        end

        169 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[32] = localMem[31] + 1;
              ip = 170;
        end

        170 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 171;
              heapClock = ~ heapClock;
        end

        171 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[577] = heapOut;                                                     // Data retrieved from heap memory
              ip = 172;
              heapClock = ~ heapClock;
        end

        172 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[33] = localMem[577];
              ip = 173;
        end

        173 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[33] == 0 ? 377 : 174;
        end

        174 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   174");
        end

        175 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   175");
        end

        176 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   176");
        end

        177 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   177");
        end

        178 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   178");
        end

        179 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   179");
        end

        180 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   180");
        end

        181 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   181");
        end

        182 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   182");
        end

        183 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   183");
        end

        184 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   184");
        end

        185 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   185");
        end

        186 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   186");
        end

        187 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   187");
        end

        188 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   188");
        end

        189 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   189");
        end

        190 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   190");
        end

        191 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   191");
        end

        192 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   192");
        end

        193 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   193");
        end

        194 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   194");
        end

        195 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   195");
        end

        196 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   196");
        end

        197 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   197");
        end

        198 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   198");
        end

        199 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   199");
        end

        200 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   200");
        end

        201 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   201");
        end

        202 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   202");
        end

        203 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   203");
        end

        204 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   204");
        end

        205 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   205");
        end

        206 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   206");
        end

        207 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   207");
        end

        208 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   208");
        end

        209 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   209");
        end

        210 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   210");
        end

        211 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   211");
        end

        212 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   212");
        end

        213 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   213");
        end

        214 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   214");
        end

        215 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   215");
        end

        216 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   216");
        end

        217 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   217");
        end

        218 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   218");
        end

        219 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   219");
        end

        220 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   220");
        end

        221 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   221");
        end

        222 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   222");
        end

        223 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   223");
        end

        224 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   224");
        end

        225 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   225");
        end

        226 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   226");
        end

        227 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   227");
        end

        228 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   228");
        end

        229 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   229");
        end

        230 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   230");
        end

        231 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   231");
        end

        232 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   232");
        end

        233 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   233");
        end

        234 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   234");
        end

        235 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   235");
        end

        236 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   236");
        end

        237 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   237");
        end

        238 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   238");
        end

        239 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   239");
        end

        240 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   240");
        end

        241 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   241");
        end

        242 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   242");
        end

        243 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   243");
        end

        244 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   244");
        end

        245 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   245");
        end

        246 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   246");
        end

        247 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   247");
        end

        248 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   248");
        end

        249 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   249");
        end

        250 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   250");
        end

        251 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   251");
        end

        252 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   252");
        end

        253 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   253");
        end

        254 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   254");
        end

        255 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   255");
        end

        256 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   256");
        end

        257 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   257");
        end

        258 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   258");
        end

        259 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   259");
        end

        260 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   260");
        end

        261 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   261");
        end

        262 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   262");
        end

        263 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   263");
        end

        264 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   264");
        end

        265 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   265");
        end

        266 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   266");
        end

        267 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   267");
        end

        268 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   268");
        end

        269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   269");
        end

        270 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   270");
        end

        271 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   271");
        end

        272 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   272");
        end

        273 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   273");
        end

        274 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   274");
        end

        275 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   275");
        end

        276 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   276");
        end

        277 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   277");
        end

        278 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   278");
        end

        279 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   279");
        end

        280 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   280");
        end

        281 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   281");
        end

        282 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   282");
        end

        283 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   283");
        end

        284 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   284");
        end

        285 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   285");
        end

        286 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   286");
        end

        287 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   287");
        end

        288 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   288");
        end

        289 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   289");
        end

        290 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   290");
        end

        291 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   291");
        end

        292 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   292");
        end

        293 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   293");
        end

        294 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   294");
        end

        295 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   295");
        end

        296 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   296");
        end

        297 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   297");
        end

        298 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   298");
        end

        299 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   299");
        end

        300 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   300");
        end

        301 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   301");
        end

        302 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   302");
        end

        303 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   303");
        end

        304 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   304");
        end

        305 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   305");
        end

        306 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   306");
        end

        307 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   307");
        end

        308 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   308");
        end

        309 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   309");
        end

        310 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   310");
        end

        311 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   311");
        end

        312 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   312");
        end

        313 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   313");
        end

        314 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   314");
        end

        315 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   315");
        end

        316 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   316");
        end

        317 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   317");
        end

        318 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   318");
        end

        319 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   319");
        end

        320 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   320");
        end

        321 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   321");
        end

        322 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   322");
        end

        323 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   323");
        end

        324 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   324");
        end

        325 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   325");
        end

        326 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   326");
        end

        327 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   327");
        end

        328 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   328");
        end

        329 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   329");
        end

        330 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   330");
        end

        331 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   331");
        end

        332 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   332");
        end

        333 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   333");
        end

        334 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   334");
        end

        335 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   335");
        end

        336 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   336");
        end

        337 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   337");
        end

        338 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   338");
        end

        339 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   339");
        end

        340 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   340");
        end

        341 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   341");
        end

        342 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   342");
        end

        343 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   343");
        end

        344 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   344");
        end

        345 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   345");
        end

        346 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   346");
        end

        347 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   347");
        end

        348 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   348");
        end

        349 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   349");
        end

        350 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   350");
        end

        351 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   351");
        end

        352 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   352");
        end

        353 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   353");
        end

        354 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   354");
        end

        355 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   355");
        end

        356 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   356");
        end

        357 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   357");
        end

        358 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   358");
        end

        359 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   359");
        end

        360 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   360");
        end

        361 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   361");
        end

        362 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   362");
        end

        363 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   363");
        end

        364 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   364");
        end

        365 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   365");
        end

        366 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   366");
        end

        367 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   367");
        end

        368 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   368");
        end

        369 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   369");
        end

        370 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   370");
        end

        371 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   371");
        end

        372 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   372");
        end

        373 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   373");
        end

        374 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   374");
        end

        375 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   375");
        end

        376 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   376");
        end

        377 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 378;
        end

        378 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 379;
              heapClock = ~ heapClock;
        end

        379 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[81] = heapOut;
              ip = 380;
        end

        380 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[635] = localMem[31];
              ip = 381;
        end

        381 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[635];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 382;
              heapClock = ~ heapClock;
        end

        382 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[636] = 0;
              ip = 383;
        end

        383 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[636];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 384;
              heapClock = ~ heapClock;
        end

        384 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 385;
              heapClock = ~ heapClock;
        end

        385 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[82] = heapOut;
              ip = 386;
        end

        386 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[637] = localMem[82];
              ip = 387;
        end

        387 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[637];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 388;
              heapClock = ~ heapClock;
        end

        388 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 389;
              heapClock = ~ heapClock;
        end

        389 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[83] = heapOut;
              ip = 390;
        end

        390 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[638] = localMem[83];
              ip = 391;
        end

        391 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[638];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 392;
              heapClock = ~ heapClock;
        end

        392 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[639] = 0;
              ip = 393;
        end

        393 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[639];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 394;
              heapClock = ~ heapClock;
        end

        394 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[640] = localMem[29];
              ip = 395;
        end

        395 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[640];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 396;
              heapClock = ~ heapClock;
        end

        396 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 397;
              heapClock = ~ heapClock;
        end

        397 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[641] = heapOut;                                                     // Data retrieved from heap memory
              ip = 398;
              heapClock = ~ heapClock;
        end

        398 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[642] = localMem[641] + 1;
              ip = 399;
        end

        399 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[29];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[642];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 400;
              heapClock = ~ heapClock;
        end

        400 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 401;
              heapClock = ~ heapClock;
        end

        401 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[643] = heapOut;                                                     // Data retrieved from heap memory
              ip = 402;
              heapClock = ~ heapClock;
        end

        402 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[644] = localMem[643];
              ip = 403;
        end

        403 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[644];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 404;
              heapClock = ~ heapClock;
        end

        404 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 405;
              heapClock = ~ heapClock;
        end

        405 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[84] = heapOut;
              ip = 406;
        end

        406 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[645] = localMem[31];
              ip = 407;
        end

        407 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[645];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 408;
              heapClock = ~ heapClock;
        end

        408 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[646] = 0;
              ip = 409;
        end

        409 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[646];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 410;
              heapClock = ~ heapClock;
        end

        410 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 411;
              heapClock = ~ heapClock;
        end

        411 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[85] = heapOut;
              ip = 412;
        end

        412 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[647] = localMem[85];
              ip = 413;
        end

        413 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[647];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 414;
              heapClock = ~ heapClock;
        end

        414 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 415;
              heapClock = ~ heapClock;
        end

        415 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[86] = heapOut;
              ip = 416;
        end

        416 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[648] = localMem[86];
              ip = 417;
        end

        417 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[648];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 418;
              heapClock = ~ heapClock;
        end

        418 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[649] = 0;
              ip = 419;
        end

        419 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[649];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 420;
              heapClock = ~ heapClock;
        end

        420 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[650] = localMem[29];
              ip = 421;
        end

        421 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[650];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 422;
              heapClock = ~ heapClock;
        end

        422 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 423;
              heapClock = ~ heapClock;
        end

        423 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[651] = heapOut;                                                     // Data retrieved from heap memory
              ip = 424;
              heapClock = ~ heapClock;
        end

        424 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[652] = localMem[651] + 1;
              ip = 425;
        end

        425 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[29];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[652];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 426;
              heapClock = ~ heapClock;
        end

        426 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 427;
              heapClock = ~ heapClock;
        end

        427 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[653] = heapOut;                                                     // Data retrieved from heap memory
              ip = 428;
              heapClock = ~ heapClock;
        end

        428 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[654] = localMem[653];
              ip = 429;
        end

        429 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[654];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 430;
              heapClock = ~ heapClock;
        end

        430 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 431;
              heapClock = ~ heapClock;
        end

        431 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[655] = heapOut;                                                     // Data retrieved from heap memory
              ip = 432;
              heapClock = ~ heapClock;
        end

        432 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[87] = !localMem[655];
              ip = 433;
        end

        433 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[87] != 0 ? 533 : 434;
        end

        434 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 435;
              heapClock = ~ heapClock;
        end

        435 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[88] = heapOut;
              ip = 436;
        end

        436 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[656] = localMem[88];
              ip = 437;
        end

        437 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[656];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 438;
              heapClock = ~ heapClock;
        end

        438 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 439;
              heapClock = ~ heapClock;
        end

        439 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[89] = heapOut;
              ip = 440;
        end

        440 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[657] = localMem[89];
              ip = 441;
        end

        441 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[657];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 442;
              heapClock = ~ heapClock;
        end

        442 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 443;
              heapClock = ~ heapClock;
        end

        443 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[658] = heapOut;                                                     // Data retrieved from heap memory
              ip = 444;
              heapClock = ~ heapClock;
        end

        444 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[90] = localMem[658];
              ip = 445;
        end

        445 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 446;
              heapClock = ~ heapClock;
        end

        446 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[659] = heapOut;                                                     // Data retrieved from heap memory
              ip = 447;
              heapClock = ~ heapClock;
        end

        447 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[91] = localMem[659];
              ip = 448;
        end

        448 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[90];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 449;
              heapClock = ~ heapClock;
        end

        449 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[91];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 450;
              heapClock = ~ heapClock;
        end

        450 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 451;
              heapClock = ~ heapClock;
        end

        451 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[660] = heapOut;                                                     // Data retrieved from heap memory
              ip = 452;
              heapClock = ~ heapClock;
        end

        452 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[92] = localMem[660];
              ip = 453;
        end

        453 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 454;
              heapClock = ~ heapClock;
        end

        454 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[661] = heapOut;                                                     // Data retrieved from heap memory
              ip = 455;
              heapClock = ~ heapClock;
        end

        455 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[93] = localMem[661];
              ip = 456;
        end

        456 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[92];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 457;
              heapClock = ~ heapClock;
        end

        457 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[93];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 458;
              heapClock = ~ heapClock;
        end

        458 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 459;
              heapClock = ~ heapClock;
        end

        459 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[662] = heapOut;                                                     // Data retrieved from heap memory
              ip = 460;
              heapClock = ~ heapClock;
        end

        460 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[94] = localMem[662];
              ip = 461;
        end

        461 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 462;
              heapClock = ~ heapClock;
        end

        462 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[663] = heapOut;                                                     // Data retrieved from heap memory
              ip = 463;
              heapClock = ~ heapClock;
        end

        463 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[95] = localMem[663];
              ip = 464;
        end

        464 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[96] = localMem[31] + 1;
              ip = 465;
        end

        465 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[94];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 466;
              heapClock = ~ heapClock;
        end

        466 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[95];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[96];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 467;
              heapClock = ~ heapClock;
        end

        467 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 468;
              heapClock = ~ heapClock;
        end

        468 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[664] = heapOut;                                                     // Data retrieved from heap memory
              ip = 469;
              heapClock = ~ heapClock;
        end

        469 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[97] = localMem[664];
              ip = 470;
        end

        470 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 471;
              heapClock = ~ heapClock;
        end

        471 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[665] = heapOut;                                                     // Data retrieved from heap memory
              ip = 472;
              heapClock = ~ heapClock;
        end

        472 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[98] = localMem[665];
              ip = 473;
        end

        473 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[97];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 474;
              heapClock = ~ heapClock;
        end

        474 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[98];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 475;
              heapClock = ~ heapClock;
        end

        475 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 476;
              heapClock = ~ heapClock;
        end

        476 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[666] = heapOut;                                                     // Data retrieved from heap memory
              ip = 477;
              heapClock = ~ heapClock;
        end

        477 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[99] = localMem[666];
              ip = 478;
        end

        478 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 479;
              heapClock = ~ heapClock;
        end

        479 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[667] = heapOut;                                                     // Data retrieved from heap memory
              ip = 480;
              heapClock = ~ heapClock;
        end

        480 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[100] = localMem[667];
              ip = 481;
        end

        481 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[99];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 482;
              heapClock = ~ heapClock;
        end

        482 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[100];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 483;
              heapClock = ~ heapClock;
        end

        483 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 484;
              heapClock = ~ heapClock;
        end

        484 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[668] = heapOut;                                                     // Data retrieved from heap memory
              ip = 485;
              heapClock = ~ heapClock;
        end

        485 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[101] = localMem[668];
              ip = 486;
        end

        486 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 487;
              heapClock = ~ heapClock;
        end

        487 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[669] = heapOut;                                                     // Data retrieved from heap memory
              ip = 488;
              heapClock = ~ heapClock;
        end

        488 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[102] = localMem[669];
              ip = 489;
        end

        489 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[103] = localMem[31] + 1;
              ip = 490;
        end

        490 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[101];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 491;
              heapClock = ~ heapClock;
        end

        491 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[102];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[103];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 492;
              heapClock = ~ heapClock;
        end

        492 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 493;
              heapClock = ~ heapClock;
        end

        493 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[670] = heapOut;                                                     // Data retrieved from heap memory
              ip = 494;
              heapClock = ~ heapClock;
        end

        494 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[104] = localMem[670];
              ip = 495;
        end

        495 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[105] = localMem[104] + 1;
              ip = 496;
        end

        496 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 497;
              heapClock = ~ heapClock;
        end

        497 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[671] = heapOut;                                                     // Data retrieved from heap memory
              ip = 498;
              heapClock = ~ heapClock;
        end

        498 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[106] = localMem[671];
              ip = 499;
        end

        499 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 500;
        end

        500 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[107] = 0;
              ip = 501;
        end

        501 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 502;
        end

        502 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[107] >= localMem[105] ? 511 : 503;
        end

        503 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[106];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[107];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 504;
              heapClock = ~ heapClock;
        end

        504 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[672] = heapOut;                                                     // Data retrieved from heap memory
              ip = 505;
              heapClock = ~ heapClock;
        end

        505 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[108] = localMem[672];
              ip = 506;
        end

        506 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[673] = localMem[81];
              ip = 507;
        end

        507 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[108];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[673];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 508;
              heapClock = ~ heapClock;
        end

        508 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 509;
        end

        509 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[107] = localMem[107] + 1;
              ip = 510;
        end

        510 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 501;
        end

        511 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 512;
        end

        512 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 513;
              heapClock = ~ heapClock;
        end

        513 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[674] = heapOut;                                                     // Data retrieved from heap memory
              ip = 514;
              heapClock = ~ heapClock;
        end

        514 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[109] = localMem[674];
              ip = 515;
        end

        515 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[110] = localMem[109] + 1;
              ip = 516;
        end

        516 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 517;
              heapClock = ~ heapClock;
        end

        517 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[675] = heapOut;                                                     // Data retrieved from heap memory
              ip = 518;
              heapClock = ~ heapClock;
        end

        518 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[111] = localMem[675];
              ip = 519;
        end

        519 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 520;
        end

        520 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[112] = 0;
              ip = 521;
        end

        521 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 522;
        end

        522 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[112] >= localMem[110] ? 531 : 523;
        end

        523 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[111];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[112];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 524;
              heapClock = ~ heapClock;
        end

        524 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[676] = heapOut;                                                     // Data retrieved from heap memory
              ip = 525;
              heapClock = ~ heapClock;
        end

        525 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[113] = localMem[676];
              ip = 526;
        end

        526 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[677] = localMem[84];
              ip = 527;
        end

        527 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[113];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[677];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 528;
              heapClock = ~ heapClock;
        end

        528 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 529;
        end

        529 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[112] = localMem[112] + 1;
              ip = 530;
        end

        530 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 521;
        end

        531 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 532;
        end

        532 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 570;
        end

        533 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 534;
        end

        534 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 535;
              heapClock = ~ heapClock;
        end

        535 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[114] = heapOut;
              ip = 536;
        end

        536 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[678] = localMem[114];
              ip = 537;
        end

        537 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[26];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[678];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 538;
              heapClock = ~ heapClock;
        end

        538 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 539;
              heapClock = ~ heapClock;
        end

        539 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[679] = heapOut;                                                     // Data retrieved from heap memory
              ip = 540;
              heapClock = ~ heapClock;
        end

        540 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[115] = localMem[679];
              ip = 541;
        end

        541 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 542;
              heapClock = ~ heapClock;
        end

        542 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[680] = heapOut;                                                     // Data retrieved from heap memory
              ip = 543;
              heapClock = ~ heapClock;
        end

        543 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[116] = localMem[680];
              ip = 544;
        end

        544 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[115];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 545;
              heapClock = ~ heapClock;
        end

        545 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[116];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 546;
              heapClock = ~ heapClock;
        end

        546 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 547;
              heapClock = ~ heapClock;
        end

        547 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[681] = heapOut;                                                     // Data retrieved from heap memory
              ip = 548;
              heapClock = ~ heapClock;
        end

        548 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[117] = localMem[681];
              ip = 549;
        end

        549 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 550;
              heapClock = ~ heapClock;
        end

        550 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[682] = heapOut;                                                     // Data retrieved from heap memory
              ip = 551;
              heapClock = ~ heapClock;
        end

        551 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[118] = localMem[682];
              ip = 552;
        end

        552 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[117];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 553;
              heapClock = ~ heapClock;
        end

        553 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[118];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 554;
              heapClock = ~ heapClock;
        end

        554 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 555;
              heapClock = ~ heapClock;
        end

        555 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[683] = heapOut;                                                     // Data retrieved from heap memory
              ip = 556;
              heapClock = ~ heapClock;
        end

        556 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[119] = localMem[683];
              ip = 557;
        end

        557 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 558;
              heapClock = ~ heapClock;
        end

        558 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[684] = heapOut;                                                     // Data retrieved from heap memory
              ip = 559;
              heapClock = ~ heapClock;
        end

        559 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[120] = localMem[684];
              ip = 560;
        end

        560 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[119];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 561;
              heapClock = ~ heapClock;
        end

        561 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[120];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 562;
              heapClock = ~ heapClock;
        end

        562 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 563;
              heapClock = ~ heapClock;
        end

        563 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[685] = heapOut;                                                     // Data retrieved from heap memory
              ip = 564;
              heapClock = ~ heapClock;
        end

        564 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[121] = localMem[685];
              ip = 565;
        end

        565 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 566;
              heapClock = ~ heapClock;
        end

        566 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[686] = heapOut;                                                     // Data retrieved from heap memory
              ip = 567;
              heapClock = ~ heapClock;
        end

        567 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[122] = localMem[686];
              ip = 568;
        end

        568 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[121];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 569;
              heapClock = ~ heapClock;
        end

        569 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[122];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 570;
              heapClock = ~ heapClock;
        end

        570 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 571;
        end

        571 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[687] = localMem[26];
              ip = 572;
        end

        572 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[687];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 573;
              heapClock = ~ heapClock;
        end

        573 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[688] = localMem[26];
              ip = 574;
        end

        574 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[688];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 575;
              heapClock = ~ heapClock;
        end

        575 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 576;
              heapClock = ~ heapClock;
        end

        576 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[689] = heapOut;                                                     // Data retrieved from heap memory
              ip = 577;
              heapClock = ~ heapClock;
        end

        577 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[123] = localMem[689];
              ip = 578;
        end

        578 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[123];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 579;
              heapClock = ~ heapClock;
        end

        579 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[690] = heapOut;                                                     // Data retrieved from heap memory
              ip = 580;
              heapClock = ~ heapClock;
        end

        580 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[124] = localMem[690];
              ip = 581;
        end

        581 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 582;
              heapClock = ~ heapClock;
        end

        582 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[691] = heapOut;                                                     // Data retrieved from heap memory
              ip = 583;
              heapClock = ~ heapClock;
        end

        583 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[125] = localMem[691];
              ip = 584;
        end

        584 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[125];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 585;
              heapClock = ~ heapClock;
        end

        585 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[692] = heapOut;                                                     // Data retrieved from heap memory
              ip = 586;
              heapClock = ~ heapClock;
        end

        586 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[126] = localMem[692];
              ip = 587;
        end

        587 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 588;
              heapClock = ~ heapClock;
        end

        588 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[693] = heapOut;                                                     // Data retrieved from heap memory
              ip = 589;
              heapClock = ~ heapClock;
        end

        589 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[127] = localMem[693];
              ip = 590;
        end

        590 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[694] = localMem[124];
              ip = 591;
        end

        591 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[127];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[694];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 592;
              heapClock = ~ heapClock;
        end

        592 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 593;
              heapClock = ~ heapClock;
        end

        593 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[695] = heapOut;                                                     // Data retrieved from heap memory
              ip = 594;
              heapClock = ~ heapClock;
        end

        594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[128] = localMem[695];
              ip = 595;
        end

        595 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[696] = localMem[126];
              ip = 596;
        end

        596 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[128];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[696];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 597;
              heapClock = ~ heapClock;
        end

        597 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 598;
              heapClock = ~ heapClock;
        end

        598 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[697] = heapOut;                                                     // Data retrieved from heap memory
              ip = 599;
              heapClock = ~ heapClock;
        end

        599 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[129] = localMem[697];
              ip = 600;
        end

        600 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[698] = localMem[81];
              ip = 601;
        end

        601 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[129];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[698];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 602;
              heapClock = ~ heapClock;
        end

        602 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 603;
              heapClock = ~ heapClock;
        end

        603 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[699] = heapOut;                                                     // Data retrieved from heap memory
              ip = 604;
              heapClock = ~ heapClock;
        end

        604 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[130] = localMem[699];
              ip = 605;
        end

        605 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[700] = localMem[84];
              ip = 606;
        end

        606 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[130];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[700];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 607;
              heapClock = ~ heapClock;
        end

        607 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[701] = 1;
              ip = 608;
        end

        608 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[26];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[701];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 609;
              heapClock = ~ heapClock;
        end

        609 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 610;
              heapClock = ~ heapClock;
        end

        610 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[702] = heapOut;                                                     // Data retrieved from heap memory
              ip = 611;
              heapClock = ~ heapClock;
        end

        611 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[131] = localMem[702];
              ip = 612;
        end

        612 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[131];
              ip = 613;
              heapClock = ~ heapClock;
        end

        613 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 614;
              heapClock = ~ heapClock;
        end

        614 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[703] = heapOut;                                                     // Data retrieved from heap memory
              ip = 615;
              heapClock = ~ heapClock;
        end

        615 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[132] = localMem[703];
              ip = 616;
        end

        616 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[132];
              ip = 617;
              heapClock = ~ heapClock;
        end

        617 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 618;
              heapClock = ~ heapClock;
        end

        618 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[704] = heapOut;                                                     // Data retrieved from heap memory
              ip = 619;
              heapClock = ~ heapClock;
        end

        619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[133] = localMem[704];
              ip = 620;
        end

        620 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 2;
              heapArray  = localMem[133];
              ip = 621;
              heapClock = ~ heapClock;
        end

        621 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 623;
        end

        622 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   622");
        end

        623 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 624;
        end

        624 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[27] = 1;
              ip = 625;
        end

        625 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 628;
        end

        626 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 627;
        end

        627 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[27] = 0;
              ip = 628;
        end

        628 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 629;
        end

        629 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 630;
        end

        630 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 631;
        end

        631 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[134] = 0;
              ip = 632;
        end

        632 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 633;
        end

        633 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[134] >= 99 ? 1654 : 634;
        end

        634 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 635;
              heapClock = ~ heapClock;
        end

        635 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[705] = heapOut;                                                     // Data retrieved from heap memory
              ip = 636;
              heapClock = ~ heapClock;
        end

        636 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[135] = localMem[705];
              ip = 637;
        end

        637 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[136] = localMem[135] - 1;
              ip = 638;
        end

        638 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 639;
              heapClock = ~ heapClock;
        end

        639 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[706] = heapOut;                                                     // Data retrieved from heap memory
              ip = 640;
              heapClock = ~ heapClock;
        end

        640 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[137] = localMem[706];
              ip = 641;
        end

        641 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[137];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[136];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 642;
              heapClock = ~ heapClock;
        end

        642 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[707] = heapOut;                                                     // Data retrieved from heap memory
              ip = 643;
              heapClock = ~ heapClock;
        end

        643 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[138] = localMem[707];
              ip = 644;
        end

        644 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[1] <= localMem[138] ? 1140 : 645;
        end

        645 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 646;
              heapClock = ~ heapClock;
        end

        646 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[708] = heapOut;                                                     // Data retrieved from heap memory
              ip = 647;
              heapClock = ~ heapClock;
        end

        647 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[139] = !localMem[708];
              ip = 648;
        end

        648 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[139] == 0 ? 656 : 649;
        end

        649 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[709] = localMem[26];
              ip = 650;
        end

        650 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[709];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 651;
              heapClock = ~ heapClock;
        end

        651 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[710] = 2;
              ip = 652;
        end

        652 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[710];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 653;
              heapClock = ~ heapClock;
        end

        653 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[711] = localMem[135] - 1;
              ip = 654;
        end

        654 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[711];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 655;
              heapClock = ~ heapClock;
        end

        655 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1658;
        end

        656 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 657;
        end

        657 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 658;
              heapClock = ~ heapClock;
        end

        658 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[712] = heapOut;                                                     // Data retrieved from heap memory
              ip = 659;
              heapClock = ~ heapClock;
        end

        659 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[140] = localMem[712];
              ip = 660;
        end

        660 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[135];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 661;
              heapClock = ~ heapClock;
        end

        661 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[713] = heapOut;                                                     // Data retrieved from heap memory
              ip = 662;
              heapClock = ~ heapClock;
        end

        662 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[141] = localMem[713];
              ip = 663;
        end

        663 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 664;
        end

        664 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 665;
              heapClock = ~ heapClock;
        end

        665 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[714] = heapOut;                                                     // Data retrieved from heap memory
              ip = 666;
              heapClock = ~ heapClock;
        end

        666 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[143] = localMem[714];
              ip = 667;
        end

        667 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 668;
              heapClock = ~ heapClock;
        end

        668 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[715] = heapOut;                                                     // Data retrieved from heap memory
              ip = 669;
              heapClock = ~ heapClock;
        end

        669 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[144] = localMem[715];
              ip = 670;
        end

        670 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 671;
              heapClock = ~ heapClock;
        end

        671 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[716] = heapOut;                                                     // Data retrieved from heap memory
              ip = 672;
              heapClock = ~ heapClock;
        end

        672 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[145] = localMem[716];
              ip = 673;
        end

        673 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[143] <  localMem[145] ? 1133 : 674;
        end

        674 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[146] = localMem[145];
              ip = 675;
        end

        675 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[146] = localMem[146] >> 1;
              ip = 676;
              ip = 676;
        end

        676 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[147] = localMem[146] + 1;
              ip = 677;
        end

        677 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 678;
              heapClock = ~ heapClock;
        end

        678 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[717] = heapOut;                                                     // Data retrieved from heap memory
              ip = 679;
              heapClock = ~ heapClock;
        end

        679 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[148] = localMem[717];
              ip = 680;
        end

        680 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[148] == 0 ? 884 : 681;
        end

        681 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 682;
              heapClock = ~ heapClock;
        end

        682 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[149] = heapOut;
              ip = 683;
        end

        683 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[718] = localMem[146];
              ip = 684;
        end

        684 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[718];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 685;
              heapClock = ~ heapClock;
        end

        685 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[719] = 0;
              ip = 686;
        end

        686 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[719];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 687;
              heapClock = ~ heapClock;
        end

        687 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 688;
              heapClock = ~ heapClock;
        end

        688 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[150] = heapOut;
              ip = 689;
        end

        689 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[720] = localMem[150];
              ip = 690;
        end

        690 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[720];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 691;
              heapClock = ~ heapClock;
        end

        691 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 692;
              heapClock = ~ heapClock;
        end

        692 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[151] = heapOut;
              ip = 693;
        end

        693 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[721] = localMem[151];
              ip = 694;
        end

        694 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[721];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 695;
              heapClock = ~ heapClock;
        end

        695 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[722] = 0;
              ip = 696;
        end

        696 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[722];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 697;
              heapClock = ~ heapClock;
        end

        697 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[723] = localMem[144];
              ip = 698;
        end

        698 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[723];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 699;
              heapClock = ~ heapClock;
        end

        699 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 700;
              heapClock = ~ heapClock;
        end

        700 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[724] = heapOut;                                                     // Data retrieved from heap memory
              ip = 701;
              heapClock = ~ heapClock;
        end

        701 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[725] = localMem[724] + 1;
              ip = 702;
        end

        702 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[144];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[725];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 703;
              heapClock = ~ heapClock;
        end

        703 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 704;
              heapClock = ~ heapClock;
        end

        704 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[726] = heapOut;                                                     // Data retrieved from heap memory
              ip = 705;
              heapClock = ~ heapClock;
        end

        705 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[727] = localMem[726];
              ip = 706;
        end

        706 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[727];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 707;
              heapClock = ~ heapClock;
        end

        707 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 708;
              heapClock = ~ heapClock;
        end

        708 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[728] = heapOut;                                                     // Data retrieved from heap memory
              ip = 709;
              heapClock = ~ heapClock;
        end

        709 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[152] = !localMem[728];
              ip = 710;
        end

        710 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[152] != 0 ? 765 : 711;
        end

        711 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 712;
              heapClock = ~ heapClock;
        end

        712 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[153] = heapOut;
              ip = 713;
        end

        713 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[729] = localMem[153];
              ip = 714;
        end

        714 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[729];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 715;
              heapClock = ~ heapClock;
        end

        715 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 716;
              heapClock = ~ heapClock;
        end

        716 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[730] = heapOut;                                                     // Data retrieved from heap memory
              ip = 717;
              heapClock = ~ heapClock;
        end

        717 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[154] = localMem[730];
              ip = 718;
        end

        718 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 719;
              heapClock = ~ heapClock;
        end

        719 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[731] = heapOut;                                                     // Data retrieved from heap memory
              ip = 720;
              heapClock = ~ heapClock;
        end

        720 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[155] = localMem[731];
              ip = 721;
        end

        721 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[154];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 722;
              heapClock = ~ heapClock;
        end

        722 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[155];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[146];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 723;
              heapClock = ~ heapClock;
        end

        723 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 724;
              heapClock = ~ heapClock;
        end

        724 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[732] = heapOut;                                                     // Data retrieved from heap memory
              ip = 725;
              heapClock = ~ heapClock;
        end

        725 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[156] = localMem[732];
              ip = 726;
        end

        726 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 727;
              heapClock = ~ heapClock;
        end

        727 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[733] = heapOut;                                                     // Data retrieved from heap memory
              ip = 728;
              heapClock = ~ heapClock;
        end

        728 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[157] = localMem[733];
              ip = 729;
        end

        729 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[156];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 730;
              heapClock = ~ heapClock;
        end

        730 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[157];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[146];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 731;
              heapClock = ~ heapClock;
        end

        731 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 732;
              heapClock = ~ heapClock;
        end

        732 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[734] = heapOut;                                                     // Data retrieved from heap memory
              ip = 733;
              heapClock = ~ heapClock;
        end

        733 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[158] = localMem[734];
              ip = 734;
        end

        734 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 735;
              heapClock = ~ heapClock;
        end

        735 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[735] = heapOut;                                                     // Data retrieved from heap memory
              ip = 736;
              heapClock = ~ heapClock;
        end

        736 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[159] = localMem[735];
              ip = 737;
        end

        737 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[160] = localMem[146] + 1;
              ip = 738;
        end

        738 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[158];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 739;
              heapClock = ~ heapClock;
        end

        739 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[159];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[160];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 740;
              heapClock = ~ heapClock;
        end

        740 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 741;
              heapClock = ~ heapClock;
        end

        741 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[736] = heapOut;                                                     // Data retrieved from heap memory
              ip = 742;
              heapClock = ~ heapClock;
        end

        742 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[161] = localMem[736];
              ip = 743;
        end

        743 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[162] = localMem[161] + 1;
              ip = 744;
        end

        744 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 745;
              heapClock = ~ heapClock;
        end

        745 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[737] = heapOut;                                                     // Data retrieved from heap memory
              ip = 746;
              heapClock = ~ heapClock;
        end

        746 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[163] = localMem[737];
              ip = 747;
        end

        747 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 748;
        end

        748 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[164] = 0;
              ip = 749;
        end

        749 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 750;
        end

        750 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[164] >= localMem[162] ? 759 : 751;
        end

        751 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[163];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[164];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 752;
              heapClock = ~ heapClock;
        end

        752 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[738] = heapOut;                                                     // Data retrieved from heap memory
              ip = 753;
              heapClock = ~ heapClock;
        end

        753 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[165] = localMem[738];
              ip = 754;
        end

        754 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[739] = localMem[149];
              ip = 755;
        end

        755 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[165];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[739];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 756;
              heapClock = ~ heapClock;
        end

        756 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 757;
        end

        757 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[164] = localMem[164] + 1;
              ip = 758;
        end

        758 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 749;
        end

        759 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 760;
        end

        760 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 761;
              heapClock = ~ heapClock;
        end

        761 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[740] = heapOut;                                                     // Data retrieved from heap memory
              ip = 762;
              heapClock = ~ heapClock;
        end

        762 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[166] = localMem[740];
              ip = 763;
        end

        763 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[147];
              heapArray  = localMem[166];
              ip = 764;
              heapClock = ~ heapClock;
        end

        764 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 782;
        end

        765 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   765");
        end

        766 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   766");
        end

        767 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   767");
        end

        768 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   768");
        end

        769 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   769");
        end

        770 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   770");
        end

        771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   771");
        end

        772 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   772");
        end

        773 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   773");
        end

        774 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   774");
        end

        775 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   775");
        end

        776 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   776");
        end

        777 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   777");
        end

        778 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   778");
        end

        779 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   779");
        end

        780 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   780");
        end

        781 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   781");
        end

        782 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 783;
        end

        783 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[745] = localMem[146];
              ip = 784;
        end

        784 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[141];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[745];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 785;
              heapClock = ~ heapClock;
        end

        785 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[746] = localMem[148];
              ip = 786;
        end

        786 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[746];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 787;
              heapClock = ~ heapClock;
        end

        787 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 788;
              heapClock = ~ heapClock;
        end

        788 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[747] = heapOut;                                                     // Data retrieved from heap memory
              ip = 789;
              heapClock = ~ heapClock;
        end

        789 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[171] = localMem[747];
              ip = 790;
        end

        790 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 791;
              heapClock = ~ heapClock;
        end

        791 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[748] = heapOut;                                                     // Data retrieved from heap memory
              ip = 792;
              heapClock = ~ heapClock;
        end

        792 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[172] = localMem[748];
              ip = 793;
        end

        793 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[172];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[171];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 794;
              heapClock = ~ heapClock;
        end

        794 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[749] = heapOut;                                                     // Data retrieved from heap memory
              ip = 795;
              heapClock = ~ heapClock;
        end

        795 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[173] = localMem[749];
              ip = 796;
        end

        796 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[173] != localMem[141] ? 837 : 797;
        end

        797 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 798;
              heapClock = ~ heapClock;
        end

        798 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[750] = heapOut;                                                     // Data retrieved from heap memory
              ip = 799;
              heapClock = ~ heapClock;
        end

        799 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[174] = localMem[750];
              ip = 800;
        end

        800 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[174];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[146];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 801;
              heapClock = ~ heapClock;
        end

        801 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[751] = heapOut;                                                     // Data retrieved from heap memory
              ip = 802;
              heapClock = ~ heapClock;
        end

        802 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[175] = localMem[751];
              ip = 803;
        end

        803 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 804;
              heapClock = ~ heapClock;
        end

        804 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[752] = heapOut;                                                     // Data retrieved from heap memory
              ip = 805;
              heapClock = ~ heapClock;
        end

        805 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[176] = localMem[752];
              ip = 806;
        end

        806 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[753] = localMem[175];
              ip = 807;
        end

        807 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[176];                                                // Array to write to
              heapIndex   = localMem[171];                                                // Index of element to write to
              heapIn      = localMem[753];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 808;
              heapClock = ~ heapClock;
        end

        808 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 809;
              heapClock = ~ heapClock;
        end

        809 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[754] = heapOut;                                                     // Data retrieved from heap memory
              ip = 810;
              heapClock = ~ heapClock;
        end

        810 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[177] = localMem[754];
              ip = 811;
        end

        811 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[177];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[146];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 812;
              heapClock = ~ heapClock;
        end

        812 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[755] = heapOut;                                                     // Data retrieved from heap memory
              ip = 813;
              heapClock = ~ heapClock;
        end

        813 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[178] = localMem[755];
              ip = 814;
        end

        814 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 815;
              heapClock = ~ heapClock;
        end

        815 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[756] = heapOut;                                                     // Data retrieved from heap memory
              ip = 816;
              heapClock = ~ heapClock;
        end

        816 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[179] = localMem[756];
              ip = 817;
        end

        817 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[757] = localMem[178];
              ip = 818;
        end

        818 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[179];                                                // Array to write to
              heapIndex   = localMem[171];                                                // Index of element to write to
              heapIn      = localMem[757];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 819;
              heapClock = ~ heapClock;
        end

        819 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 820;
              heapClock = ~ heapClock;
        end

        820 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[758] = heapOut;                                                     // Data retrieved from heap memory
              ip = 821;
              heapClock = ~ heapClock;
        end

        821 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[180] = localMem[758];
              ip = 822;
        end

        822 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[146];
              heapArray  = localMem[180];
              ip = 823;
              heapClock = ~ heapClock;
        end

        823 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 824;
              heapClock = ~ heapClock;
        end

        824 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[759] = heapOut;                                                     // Data retrieved from heap memory
              ip = 825;
              heapClock = ~ heapClock;
        end

        825 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[181] = localMem[759];
              ip = 826;
        end

        826 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[146];
              heapArray  = localMem[181];
              ip = 827;
              heapClock = ~ heapClock;
        end

        827 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[182] = localMem[171] + 1;
              ip = 828;
        end

        828 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[760] = localMem[182];
              ip = 829;
        end

        829 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[148];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[760];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 830;
              heapClock = ~ heapClock;
        end

        830 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 831;
              heapClock = ~ heapClock;
        end

        831 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[761] = heapOut;                                                     // Data retrieved from heap memory
              ip = 832;
              heapClock = ~ heapClock;
        end

        832 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[183] = localMem[761];
              ip = 833;
        end

        833 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[762] = localMem[149];
              ip = 834;
        end

        834 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[183];                                                // Array to write to
              heapIndex   = localMem[182];                                                // Index of element to write to
              heapIn      = localMem[762];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 835;
              heapClock = ~ heapClock;
        end

        835 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1130;
        end

        836 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   836");
        end

        837 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   837");
        end

        838 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   838");
        end

        839 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   839");
        end

        840 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   840");
        end

        841 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   841");
        end

        842 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   842");
        end

        843 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   843");
        end

        844 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   844");
        end

        845 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   845");
        end

        846 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   846");
        end

        847 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   847");
        end

        848 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   848");
        end

        849 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   849");
        end

        850 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   850");
        end

        851 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   851");
        end

        852 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   852");
        end

        853 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   853");
        end

        854 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   854");
        end

        855 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   855");
        end

        856 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   856");
        end

        857 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   857");
        end

        858 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   858");
        end

        859 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   859");
        end

        860 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   860");
        end

        861 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   861");
        end

        862 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   862");
        end

        863 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   863");
        end

        864 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   864");
        end

        865 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   865");
        end

        866 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   866");
        end

        867 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   867");
        end

        868 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   868");
        end

        869 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   869");
        end

        870 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   870");
        end

        871 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   871");
        end

        872 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   872");
        end

        873 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   873");
        end

        874 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   874");
        end

        875 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   875");
        end

        876 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   876");
        end

        877 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   877");
        end

        878 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   878");
        end

        879 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   879");
        end

        880 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   880");
        end

        881 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   881");
        end

        882 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   882");
        end

        883 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   883");
        end

        884 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   884");
        end

        885 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   885");
        end

        886 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   886");
        end

        887 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   887");
        end

        888 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   888");
        end

        889 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   889");
        end

        890 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   890");
        end

        891 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   891");
        end

        892 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   892");
        end

        893 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   893");
        end

        894 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   894");
        end

        895 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   895");
        end

        896 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   896");
        end

        897 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   897");
        end

        898 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   898");
        end

        899 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   899");
        end

        900 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   900");
        end

        901 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   901");
        end

        902 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   902");
        end

        903 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   903");
        end

        904 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   904");
        end

        905 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   905");
        end

        906 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   906");
        end

        907 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   907");
        end

        908 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   908");
        end

        909 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   909");
        end

        910 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   910");
        end

        911 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   911");
        end

        912 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   912");
        end

        913 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   913");
        end

        914 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   914");
        end

        915 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   915");
        end

        916 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   916");
        end

        917 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   917");
        end

        918 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   918");
        end

        919 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   919");
        end

        920 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   920");
        end

        921 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   921");
        end

        922 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   922");
        end

        923 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   923");
        end

        924 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   924");
        end

        925 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   925");
        end

        926 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   926");
        end

        927 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   927");
        end

        928 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   928");
        end

        929 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   929");
        end

        930 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   930");
        end

        931 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   931");
        end

        932 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   932");
        end

        933 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   933");
        end

        934 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   934");
        end

        935 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   935");
        end

        936 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   936");
        end

        937 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   937");
        end

        938 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   938");
        end

        939 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   939");
        end

        940 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   940");
        end

        941 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   941");
        end

        942 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   942");
        end

        943 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   943");
        end

        944 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   944");
        end

        945 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   945");
        end

        946 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   946");
        end

        947 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   947");
        end

        948 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   948");
        end

        949 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   949");
        end

        950 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   950");
        end

        951 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   951");
        end

        952 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   952");
        end

        953 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   953");
        end

        954 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   954");
        end

        955 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   955");
        end

        956 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   956");
        end

        957 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   957");
        end

        958 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   958");
        end

        959 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   959");
        end

        960 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   960");
        end

        961 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   961");
        end

        962 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   962");
        end

        963 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   963");
        end

        964 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   964");
        end

        965 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   965");
        end

        966 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   966");
        end

        967 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   967");
        end

        968 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   968");
        end

        969 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   969");
        end

        970 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   970");
        end

        971 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   971");
        end

        972 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   972");
        end

        973 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   973");
        end

        974 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   974");
        end

        975 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   975");
        end

        976 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   976");
        end

        977 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   977");
        end

        978 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   978");
        end

        979 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   979");
        end

        980 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   980");
        end

        981 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   981");
        end

        982 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   982");
        end

        983 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   983");
        end

        984 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   984");
        end

        985 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   985");
        end

        986 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   986");
        end

        987 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   987");
        end

        988 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   988");
        end

        989 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   989");
        end

        990 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   990");
        end

        991 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   991");
        end

        992 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   992");
        end

        993 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   993");
        end

        994 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   994");
        end

        995 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   995");
        end

        996 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   996");
        end

        997 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   997");
        end

        998 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   998");
        end

        999 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   999");
        end

       1000 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1000");
        end

       1001 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1001");
        end

       1002 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1002");
        end

       1003 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1003");
        end

       1004 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1004");
        end

       1005 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1005");
        end

       1006 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1006");
        end

       1007 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1007");
        end

       1008 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1008");
        end

       1009 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1009");
        end

       1010 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1010");
        end

       1011 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1011");
        end

       1012 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1012");
        end

       1013 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1013");
        end

       1014 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1014");
        end

       1015 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1015");
        end

       1016 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1016");
        end

       1017 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1017");
        end

       1018 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1018");
        end

       1019 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1019");
        end

       1020 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1020");
        end

       1021 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1021");
        end

       1022 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1022");
        end

       1023 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1023");
        end

       1024 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1024");
        end

       1025 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1025");
        end

       1026 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1026");
        end

       1027 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1027");
        end

       1028 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1028");
        end

       1029 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1029");
        end

       1030 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1030");
        end

       1031 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1031");
        end

       1032 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1032");
        end

       1033 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1033");
        end

       1034 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1034");
        end

       1035 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1035");
        end

       1036 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1036");
        end

       1037 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1037");
        end

       1038 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1038");
        end

       1039 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1039");
        end

       1040 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1040");
        end

       1041 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1041");
        end

       1042 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1042");
        end

       1043 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1043");
        end

       1044 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1044");
        end

       1045 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1045");
        end

       1046 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1046");
        end

       1047 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1047");
        end

       1048 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1048");
        end

       1049 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1049");
        end

       1050 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1050");
        end

       1051 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1051");
        end

       1052 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1052");
        end

       1053 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1053");
        end

       1054 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1054");
        end

       1055 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1055");
        end

       1056 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1056");
        end

       1057 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1057");
        end

       1058 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1058");
        end

       1059 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1059");
        end

       1060 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1060");
        end

       1061 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1061");
        end

       1062 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1062");
        end

       1063 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1063");
        end

       1064 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1064");
        end

       1065 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1065");
        end

       1066 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1066");
        end

       1067 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1067");
        end

       1068 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1068");
        end

       1069 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1069");
        end

       1070 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1070");
        end

       1071 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1071");
        end

       1072 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1072");
        end

       1073 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1073");
        end

       1074 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1074");
        end

       1075 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1075");
        end

       1076 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1076");
        end

       1077 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1077");
        end

       1078 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1078");
        end

       1079 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1079");
        end

       1080 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1080");
        end

       1081 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1081");
        end

       1082 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1082");
        end

       1083 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1083");
        end

       1084 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1084");
        end

       1085 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1085");
        end

       1086 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1086");
        end

       1087 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1087");
        end

       1088 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1088");
        end

       1089 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1089");
        end

       1090 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1090");
        end

       1091 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1091");
        end

       1092 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1092");
        end

       1093 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1093");
        end

       1094 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1094");
        end

       1095 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1095");
        end

       1096 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1096");
        end

       1097 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1097");
        end

       1098 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1098");
        end

       1099 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1099");
        end

       1100 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1100");
        end

       1101 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1101");
        end

       1102 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1102");
        end

       1103 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1103");
        end

       1104 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1104");
        end

       1105 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1105");
        end

       1106 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1106");
        end

       1107 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1107");
        end

       1108 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1108");
        end

       1109 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1109");
        end

       1110 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1110");
        end

       1111 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1111");
        end

       1112 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1112");
        end

       1113 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1113");
        end

       1114 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1114");
        end

       1115 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1115");
        end

       1116 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1116");
        end

       1117 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1117");
        end

       1118 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1118");
        end

       1119 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1119");
        end

       1120 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1120");
        end

       1121 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1121");
        end

       1122 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1122");
        end

       1123 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1123");
        end

       1124 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1124");
        end

       1125 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1125");
        end

       1126 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1126");
        end

       1127 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1127");
        end

       1128 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1128");
        end

       1129 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1129");
        end

       1130 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1131;
        end

       1131 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[142] = 1;
              ip = 1132;
        end

       1132 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1135;
        end

       1133 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1134;
        end

       1134 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[142] = 0;
              ip = 1135;
        end

       1135 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1136;
        end

       1136 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[142] != 0 ? 1138 : 1137;
        end

       1137 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[26] = localMem[141];
              ip = 1138;
        end

       1138 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1139;
        end

       1139 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1651;
        end

       1140 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1140");
        end

       1141 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1141");
        end

       1142 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1142");
        end

       1143 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1143");
        end

       1144 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1144");
        end

       1145 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1145");
        end

       1146 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1146");
        end

       1147 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1147");
        end

       1148 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1148");
        end

       1149 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1149");
        end

       1150 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1150");
        end

       1151 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1151");
        end

       1152 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1152");
        end

       1153 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1153");
        end

       1154 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1154");
        end

       1155 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed  1155");
        end

       1156 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1156");
        end

       1157 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1157");
        end

       1158 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1158");
        end

       1159 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1159");
        end

       1160 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1160");
        end

       1161 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1161");
        end

       1162 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1162");
        end

       1163 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1163");
        end

       1164 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1164");
        end

       1165 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1165");
        end

       1166 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1166");
        end

       1167 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1167");
        end

       1168 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1168");
        end

       1169 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1169");
        end

       1170 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1170");
        end

       1171 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1171");
        end

       1172 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1172");
        end

       1173 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1173");
        end

       1174 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1174");
        end

       1175 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1175");
        end

       1176 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1176");
        end

       1177 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1177");
        end

       1178 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1178");
        end

       1179 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1179");
        end

       1180 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1180");
        end

       1181 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1181");
        end

       1182 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1182");
        end

       1183 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1183");
        end

       1184 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1184");
        end

       1185 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
          // $display("Should not be executed  1185");
        end

       1186 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1186");
        end

       1187 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
          // $display("Should not be executed  1187");
        end

       1188 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1188");
        end

       1189 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1189");
        end

       1190 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1190");
        end

       1191 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1191");
        end

       1192 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1192");
        end

       1193 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1193");
        end

       1194 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1194");
        end

       1195 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1195");
        end

       1196 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1196");
        end

       1197 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1197");
        end

       1198 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1198");
        end

       1199 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1199");
        end

       1200 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1200");
        end

       1201 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1201");
        end

       1202 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1202");
        end

       1203 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1203");
        end

       1204 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1204");
        end

       1205 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1205");
        end

       1206 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1206");
        end

       1207 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1207");
        end

       1208 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1208");
        end

       1209 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1209");
        end

       1210 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1210");
        end

       1211 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1211");
        end

       1212 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1212");
        end

       1213 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1213");
        end

       1214 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1214");
        end

       1215 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1215");
        end

       1216 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1216");
        end

       1217 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1217");
        end

       1218 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1218");
        end

       1219 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1219");
        end

       1220 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1220");
        end

       1221 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1221");
        end

       1222 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1222");
        end

       1223 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1223");
        end

       1224 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1224");
        end

       1225 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1225");
        end

       1226 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1226");
        end

       1227 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1227");
        end

       1228 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1228");
        end

       1229 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1229");
        end

       1230 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1230");
        end

       1231 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1231");
        end

       1232 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1232");
        end

       1233 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1233");
        end

       1234 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1234");
        end

       1235 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1235");
        end

       1236 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1236");
        end

       1237 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1237");
        end

       1238 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1238");
        end

       1239 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1239");
        end

       1240 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1240");
        end

       1241 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1241");
        end

       1242 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1242");
        end

       1243 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1243");
        end

       1244 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1244");
        end

       1245 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1245");
        end

       1246 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1246");
        end

       1247 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1247");
        end

       1248 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1248");
        end

       1249 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1249");
        end

       1250 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1250");
        end

       1251 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1251");
        end

       1252 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1252");
        end

       1253 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1253");
        end

       1254 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1254");
        end

       1255 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1255");
        end

       1256 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1256");
        end

       1257 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1257");
        end

       1258 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1258");
        end

       1259 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1259");
        end

       1260 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1260");
        end

       1261 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1261");
        end

       1262 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1262");
        end

       1263 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1263");
        end

       1264 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1264");
        end

       1265 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1265");
        end

       1266 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1266");
        end

       1267 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1267");
        end

       1268 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1268");
        end

       1269 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1269");
        end

       1270 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1270");
        end

       1271 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1271");
        end

       1272 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1272");
        end

       1273 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1273");
        end

       1274 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1274");
        end

       1275 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1275");
        end

       1276 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1276");
        end

       1277 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1277");
        end

       1278 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1278");
        end

       1279 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1279");
        end

       1280 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1280");
        end

       1281 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1281");
        end

       1282 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1282");
        end

       1283 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1283");
        end

       1284 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1284");
        end

       1285 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1285");
        end

       1286 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1286");
        end

       1287 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1287");
        end

       1288 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1288");
        end

       1289 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1289");
        end

       1290 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1290");
        end

       1291 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1291");
        end

       1292 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1292");
        end

       1293 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1293");
        end

       1294 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1294");
        end

       1295 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1295");
        end

       1296 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1296");
        end

       1297 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1297");
        end

       1298 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1298");
        end

       1299 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1299");
        end

       1300 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1300");
        end

       1301 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1301");
        end

       1302 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1302");
        end

       1303 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1303");
        end

       1304 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1304");
        end

       1305 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1305");
        end

       1306 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1306");
        end

       1307 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1307");
        end

       1308 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1308");
        end

       1309 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1309");
        end

       1310 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1310");
        end

       1311 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1311");
        end

       1312 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1312");
        end

       1313 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1313");
        end

       1314 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1314");
        end

       1315 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1315");
        end

       1316 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1316");
        end

       1317 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1317");
        end

       1318 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1318");
        end

       1319 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1319");
        end

       1320 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1320");
        end

       1321 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1321");
        end

       1322 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1322");
        end

       1323 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1323");
        end

       1324 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1324");
        end

       1325 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1325");
        end

       1326 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1326");
        end

       1327 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1327");
        end

       1328 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1328");
        end

       1329 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1329");
        end

       1330 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1330");
        end

       1331 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1331");
        end

       1332 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1332");
        end

       1333 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1333");
        end

       1334 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1334");
        end

       1335 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1335");
        end

       1336 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1336");
        end

       1337 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1337");
        end

       1338 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1338");
        end

       1339 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1339");
        end

       1340 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1340");
        end

       1341 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1341");
        end

       1342 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1342");
        end

       1343 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1343");
        end

       1344 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1344");
        end

       1345 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1345");
        end

       1346 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1346");
        end

       1347 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1347");
        end

       1348 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1348");
        end

       1349 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1349");
        end

       1350 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  1350");
        end

       1351 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1351");
        end

       1352 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1352");
        end

       1353 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1353");
        end

       1354 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1354");
        end

       1355 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1355");
        end

       1356 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1356");
        end

       1357 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1357");
        end

       1358 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1358");
        end

       1359 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1359");
        end

       1360 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1360");
        end

       1361 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1361");
        end

       1362 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1362");
        end

       1363 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1363");
        end

       1364 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1364");
        end

       1365 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1365");
        end

       1366 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1366");
        end

       1367 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1367");
        end

       1368 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1368");
        end

       1369 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1369");
        end

       1370 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1370");
        end

       1371 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1371");
        end

       1372 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1372");
        end

       1373 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1373");
        end

       1374 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1374");
        end

       1375 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1375");
        end

       1376 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1376");
        end

       1377 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1377");
        end

       1378 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1378");
        end

       1379 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1379");
        end

       1380 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1380");
        end

       1381 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1381");
        end

       1382 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1382");
        end

       1383 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1383");
        end

       1384 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1384");
        end

       1385 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1385");
        end

       1386 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1386");
        end

       1387 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1387");
        end

       1388 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1388");
        end

       1389 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1389");
        end

       1390 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1390");
        end

       1391 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1391");
        end

       1392 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1392");
        end

       1393 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1393");
        end

       1394 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1394");
        end

       1395 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1395");
        end

       1396 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1396");
        end

       1397 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1397");
        end

       1398 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1398");
        end

       1399 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1399");
        end

       1400 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1400");
        end

       1401 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1401");
        end

       1402 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1402");
        end

       1403 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1403");
        end

       1404 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1404");
        end

       1405 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1405");
        end

       1406 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1406");
        end

       1407 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1407");
        end

       1408 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1408");
        end

       1409 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1409");
        end

       1410 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1410");
        end

       1411 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1411");
        end

       1412 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1412");
        end

       1413 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1413");
        end

       1414 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1414");
        end

       1415 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1415");
        end

       1416 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1416");
        end

       1417 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1417");
        end

       1418 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1418");
        end

       1419 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1419");
        end

       1420 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1420");
        end

       1421 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1421");
        end

       1422 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1422");
        end

       1423 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1423");
        end

       1424 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1424");
        end

       1425 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1425");
        end

       1426 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1426");
        end

       1427 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1427");
        end

       1428 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1428");
        end

       1429 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1429");
        end

       1430 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1430");
        end

       1431 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1431");
        end

       1432 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1432");
        end

       1433 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1433");
        end

       1434 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1434");
        end

       1435 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1435");
        end

       1436 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1436");
        end

       1437 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1437");
        end

       1438 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1438");
        end

       1439 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1439");
        end

       1440 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1440");
        end

       1441 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1441");
        end

       1442 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1442");
        end

       1443 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1443");
        end

       1444 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1444");
        end

       1445 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1445");
        end

       1446 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1446");
        end

       1447 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1447");
        end

       1448 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1448");
        end

       1449 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1449");
        end

       1450 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1450");
        end

       1451 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1451");
        end

       1452 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1452");
        end

       1453 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1453");
        end

       1454 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1454");
        end

       1455 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1455");
        end

       1456 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1456");
        end

       1457 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1457");
        end

       1458 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1458");
        end

       1459 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1459");
        end

       1460 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1460");
        end

       1461 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1461");
        end

       1462 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1462");
        end

       1463 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1463");
        end

       1464 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1464");
        end

       1465 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1465");
        end

       1466 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1466");
        end

       1467 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1467");
        end

       1468 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1468");
        end

       1469 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1469");
        end

       1470 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1470");
        end

       1471 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1471");
        end

       1472 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1472");
        end

       1473 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1473");
        end

       1474 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1474");
        end

       1475 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1475");
        end

       1476 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1476");
        end

       1477 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1477");
        end

       1478 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1478");
        end

       1479 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1479");
        end

       1480 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1480");
        end

       1481 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1481");
        end

       1482 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1482");
        end

       1483 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1483");
        end

       1484 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1484");
        end

       1485 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1485");
        end

       1486 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1486");
        end

       1487 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1487");
        end

       1488 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1488");
        end

       1489 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1489");
        end

       1490 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1490");
        end

       1491 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1491");
        end

       1492 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1492");
        end

       1493 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1493");
        end

       1494 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1494");
        end

       1495 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1495");
        end

       1496 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1496");
        end

       1497 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1497");
        end

       1498 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1498");
        end

       1499 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1499");
        end

       1500 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1500");
        end

       1501 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1501");
        end

       1502 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1502");
        end

       1503 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1503");
        end

       1504 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1504");
        end

       1505 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1505");
        end

       1506 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1506");
        end

       1507 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1507");
        end

       1508 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1508");
        end

       1509 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1509");
        end

       1510 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1510");
        end

       1511 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1511");
        end

       1512 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1512");
        end

       1513 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1513");
        end

       1514 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1514");
        end

       1515 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1515");
        end

       1516 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1516");
        end

       1517 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1517");
        end

       1518 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1518");
        end

       1519 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1519");
        end

       1520 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1520");
        end

       1521 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1521");
        end

       1522 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1522");
        end

       1523 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1523");
        end

       1524 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1524");
        end

       1525 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1525");
        end

       1526 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1526");
        end

       1527 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1527");
        end

       1528 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1528");
        end

       1529 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1529");
        end

       1530 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1530");
        end

       1531 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1531");
        end

       1532 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1532");
        end

       1533 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1533");
        end

       1534 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1534");
        end

       1535 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1535");
        end

       1536 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1536");
        end

       1537 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1537");
        end

       1538 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1538");
        end

       1539 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1539");
        end

       1540 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1540");
        end

       1541 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1541");
        end

       1542 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1542");
        end

       1543 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1543");
        end

       1544 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1544");
        end

       1545 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1545");
        end

       1546 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1546");
        end

       1547 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1547");
        end

       1548 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1548");
        end

       1549 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1549");
        end

       1550 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1550");
        end

       1551 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1551");
        end

       1552 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1552");
        end

       1553 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1553");
        end

       1554 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1554");
        end

       1555 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1555");
        end

       1556 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1556");
        end

       1557 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1557");
        end

       1558 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1558");
        end

       1559 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1559");
        end

       1560 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1560");
        end

       1561 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1561");
        end

       1562 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1562");
        end

       1563 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1563");
        end

       1564 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1564");
        end

       1565 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1565");
        end

       1566 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1566");
        end

       1567 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1567");
        end

       1568 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1568");
        end

       1569 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1569");
        end

       1570 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1570");
        end

       1571 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1571");
        end

       1572 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1572");
        end

       1573 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1573");
        end

       1574 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1574");
        end

       1575 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1575");
        end

       1576 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1576");
        end

       1577 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1577");
        end

       1578 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1578");
        end

       1579 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1579");
        end

       1580 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1580");
        end

       1581 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1581");
        end

       1582 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1582");
        end

       1583 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1583");
        end

       1584 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1584");
        end

       1585 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1585");
        end

       1586 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1586");
        end

       1587 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1587");
        end

       1588 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1588");
        end

       1589 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1589");
        end

       1590 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1590");
        end

       1591 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1591");
        end

       1592 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1592");
        end

       1593 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1593");
        end

       1594 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1594");
        end

       1595 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1595");
        end

       1596 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1596");
        end

       1597 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1597");
        end

       1598 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1598");
        end

       1599 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1599");
        end

       1600 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1600");
        end

       1601 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1601");
        end

       1602 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1602");
        end

       1603 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1603");
        end

       1604 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1604");
        end

       1605 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1605");
        end

       1606 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1606");
        end

       1607 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1607");
        end

       1608 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1608");
        end

       1609 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1609");
        end

       1610 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1610");
        end

       1611 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1611");
        end

       1612 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1612");
        end

       1613 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1613");
        end

       1614 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1614");
        end

       1615 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1615");
        end

       1616 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1616");
        end

       1617 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1617");
        end

       1618 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1618");
        end

       1619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1619");
        end

       1620 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1620");
        end

       1621 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1621");
        end

       1622 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1622");
        end

       1623 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1623");
        end

       1624 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1624");
        end

       1625 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1625");
        end

       1626 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1626");
        end

       1627 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1627");
        end

       1628 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1628");
        end

       1629 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1629");
        end

       1630 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1630");
        end

       1631 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1631");
        end

       1632 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1632");
        end

       1633 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1633");
        end

       1634 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1634");
        end

       1635 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1635");
        end

       1636 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1636");
        end

       1637 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1637");
        end

       1638 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1638");
        end

       1639 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1639");
        end

       1640 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1640");
        end

       1641 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1641");
        end

       1642 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1642");
        end

       1643 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1643");
        end

       1644 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1644");
        end

       1645 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1645");
        end

       1646 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1646");
        end

       1647 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1647");
        end

       1648 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1648");
        end

       1649 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1649");
        end

       1650 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1650");
        end

       1651 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1652;
        end

       1652 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[134] = localMem[134] + 1;
              ip = 1653;
        end

       1653 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 632;
        end

       1654 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1654");
        end

       1655 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  1655");
        end

       1656 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1656");
        end

       1657 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1657");
        end

       1658 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1659;
        end

       1659 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1660;
              heapClock = ~ heapClock;
        end

       1660 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[986] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1661;
              heapClock = ~ heapClock;
        end

       1661 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[362] = localMem[986];
              ip = 1662;
        end

       1662 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1663;
              heapClock = ~ heapClock;
        end

       1663 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[987] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1664;
              heapClock = ~ heapClock;
        end

       1664 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[363] = localMem[987];
              ip = 1665;
        end

       1665 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1666;
              heapClock = ~ heapClock;
        end

       1666 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[988] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1667;
              heapClock = ~ heapClock;
        end

       1667 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[364] = localMem[988];
              ip = 1668;
        end

       1668 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[363] != 1 ? 1675 : 1669;
        end

       1669 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1669");
        end

       1670 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1670");
        end

       1671 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1671");
        end

       1672 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1672");
        end

       1673 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1673");
        end

       1674 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1674");
        end

       1675 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1676;
        end

       1676 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[363] != 2 ? 1691 : 1677;
        end

       1677 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[366] = localMem[364] + 1;
              ip = 1678;
        end

       1678 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1679;
              heapClock = ~ heapClock;
        end

       1679 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[991] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1680;
              heapClock = ~ heapClock;
        end

       1680 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[367] = localMem[991];
              ip = 1681;
        end

       1681 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[1];
              heapArray  = localMem[367];
              heapIndex  = localMem[366];
              ip = 1682;
              heapClock = ~ heapClock;
        end

       1682 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1683;
              heapClock = ~ heapClock;
        end

       1683 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[992] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1684;
              heapClock = ~ heapClock;
        end

       1684 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[368] = localMem[992];
              ip = 1685;
        end

       1685 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[2];
              heapArray  = localMem[368];
              heapIndex  = localMem[366];
              ip = 1686;
              heapClock = ~ heapClock;
        end

       1686 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1687;
              heapClock = ~ heapClock;
        end

       1687 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[993] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1688;
              heapClock = ~ heapClock;
        end

       1688 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[994] = localMem[993] + 1;
              ip = 1689;
        end

       1689 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[362];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[994];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1690;
              heapClock = ~ heapClock;
        end

       1690 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1704;
        end

       1691 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1691");
        end

       1692 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1692");
        end

       1693 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1693");
        end

       1694 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1694");
        end

       1695 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1695");
        end

       1696 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1696");
        end

       1697 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1697");
        end

       1698 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1698");
        end

       1699 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1699");
        end

       1700 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1700");
        end

       1701 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1701");
        end

       1702 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1702");
        end

       1703 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1703");
        end

       1704 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1705;
        end

       1705 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1706;
              heapClock = ~ heapClock;
        end

       1706 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[999] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1707;
              heapClock = ~ heapClock;
        end

       1707 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1000] = localMem[999] + 1;
              ip = 1708;
        end

       1708 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1000];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1709;
              heapClock = ~ heapClock;
        end

       1709 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1710;
        end

       1710 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1711;
              heapClock = ~ heapClock;
        end

       1711 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1001] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1712;
              heapClock = ~ heapClock;
        end

       1712 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[372] = localMem[1001];
              ip = 1713;
        end

       1713 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1714;
              heapClock = ~ heapClock;
        end

       1714 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1002] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1715;
              heapClock = ~ heapClock;
        end

       1715 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[373] = localMem[1002];
              ip = 1716;
        end

       1716 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1717;
              heapClock = ~ heapClock;
        end

       1717 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1003] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1718;
              heapClock = ~ heapClock;
        end

       1718 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[374] = localMem[1003];
              ip = 1719;
        end

       1719 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[372] <  localMem[374] ? 2179 : 1720;
        end

       1720 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[375] = localMem[374];
              ip = 1721;
        end

       1721 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[375] = localMem[375] >> 1;
              ip = 1722;
              ip = 1722;
        end

       1722 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[376] = localMem[375] + 1;
              ip = 1723;
        end

       1723 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1724;
              heapClock = ~ heapClock;
        end

       1724 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1004] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1725;
              heapClock = ~ heapClock;
        end

       1725 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[377] = localMem[1004];
              ip = 1726;
        end

       1726 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[377] == 0 ? 1930 : 1727;
        end

       1727 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1728;
              heapClock = ~ heapClock;
        end

       1728 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[378] = heapOut;
              ip = 1729;
        end

       1729 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1005] = localMem[375];
              ip = 1730;
        end

       1730 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1005];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1731;
              heapClock = ~ heapClock;
        end

       1731 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1006] = 0;
              ip = 1732;
        end

       1732 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1006];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1733;
              heapClock = ~ heapClock;
        end

       1733 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1734;
              heapClock = ~ heapClock;
        end

       1734 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[379] = heapOut;
              ip = 1735;
        end

       1735 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1007] = localMem[379];
              ip = 1736;
        end

       1736 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[1007];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1737;
              heapClock = ~ heapClock;
        end

       1737 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1738;
              heapClock = ~ heapClock;
        end

       1738 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[380] = heapOut;
              ip = 1739;
        end

       1739 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1008] = localMem[380];
              ip = 1740;
        end

       1740 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[1008];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1741;
              heapClock = ~ heapClock;
        end

       1741 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1009] = 0;
              ip = 1742;
        end

       1742 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[1009];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1743;
              heapClock = ~ heapClock;
        end

       1743 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1010] = localMem[373];
              ip = 1744;
        end

       1744 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[1010];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1745;
              heapClock = ~ heapClock;
        end

       1745 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1746;
              heapClock = ~ heapClock;
        end

       1746 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1011] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1747;
              heapClock = ~ heapClock;
        end

       1747 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1012] = localMem[1011] + 1;
              ip = 1748;
        end

       1748 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[373];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1012];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1749;
              heapClock = ~ heapClock;
        end

       1749 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1750;
              heapClock = ~ heapClock;
        end

       1750 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1013] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1751;
              heapClock = ~ heapClock;
        end

       1751 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1014] = localMem[1013];
              ip = 1752;
        end

       1752 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1014];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1753;
              heapClock = ~ heapClock;
        end

       1753 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1754;
              heapClock = ~ heapClock;
        end

       1754 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1015] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1755;
              heapClock = ~ heapClock;
        end

       1755 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[381] = !localMem[1015];
              ip = 1756;
        end

       1756 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[381] != 0 ? 1811 : 1757;
        end

       1757 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1757");
        end

       1758 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1758");
        end

       1759 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1759");
        end

       1760 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1760");
        end

       1761 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1761");
        end

       1762 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1762");
        end

       1763 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1763");
        end

       1764 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1764");
        end

       1765 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1765");
        end

       1766 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1766");
        end

       1767 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1767");
        end

       1768 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1768");
        end

       1769 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1769");
        end

       1770 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1770");
        end

       1771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1771");
        end

       1772 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1772");
        end

       1773 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1773");
        end

       1774 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1774");
        end

       1775 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1775");
        end

       1776 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1776");
        end

       1777 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1777");
        end

       1778 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1778");
        end

       1779 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1779");
        end

       1780 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1780");
        end

       1781 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1781");
        end

       1782 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1782");
        end

       1783 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1783");
        end

       1784 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1784");
        end

       1785 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1785");
        end

       1786 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1786");
        end

       1787 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1787");
        end

       1788 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1788");
        end

       1789 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1789");
        end

       1790 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1790");
        end

       1791 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1791");
        end

       1792 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1792");
        end

       1793 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1793");
        end

       1794 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1794");
        end

       1795 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1795");
        end

       1796 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1796");
        end

       1797 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1797");
        end

       1798 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1798");
        end

       1799 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1799");
        end

       1800 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1800");
        end

       1801 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1801");
        end

       1802 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1802");
        end

       1803 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1803");
        end

       1804 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1804");
        end

       1805 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1805");
        end

       1806 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1806");
        end

       1807 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1807");
        end

       1808 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1808");
        end

       1809 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1809");
        end

       1810 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1810");
        end

       1811 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1812;
        end

       1812 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1813;
              heapClock = ~ heapClock;
        end

       1813 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1028] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1814;
              heapClock = ~ heapClock;
        end

       1814 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[396] = localMem[1028];
              ip = 1815;
        end

       1815 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[378];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1816;
              heapClock = ~ heapClock;
        end

       1816 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1029] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1817;
              heapClock = ~ heapClock;
        end

       1817 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[397] = localMem[1029];
              ip = 1818;
        end

       1818 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[396];                                                 // Array to write to
              heapIndex  = localMem[376];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1819;
              heapClock = ~ heapClock;
        end

       1819 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[397];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[375];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1820;
              heapClock = ~ heapClock;
        end

       1820 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1821;
              heapClock = ~ heapClock;
        end

       1821 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1030] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1822;
              heapClock = ~ heapClock;
        end

       1822 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[398] = localMem[1030];
              ip = 1823;
        end

       1823 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[378];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1824;
              heapClock = ~ heapClock;
        end

       1824 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1031] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1825;
              heapClock = ~ heapClock;
        end

       1825 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[399] = localMem[1031];
              ip = 1826;
        end

       1826 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[398];                                                 // Array to write to
              heapIndex  = localMem[376];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1827;
              heapClock = ~ heapClock;
        end

       1827 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[399];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[375];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1828;
              heapClock = ~ heapClock;
        end

       1828 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1829;
        end

       1829 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1032] = localMem[375];
              ip = 1830;
        end

       1830 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[362];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1032];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1831;
              heapClock = ~ heapClock;
        end

       1831 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1033] = localMem[377];
              ip = 1832;
        end

       1832 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1033];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1833;
              heapClock = ~ heapClock;
        end

       1833 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1834;
              heapClock = ~ heapClock;
        end

       1834 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1034] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1835;
              heapClock = ~ heapClock;
        end

       1835 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[400] = localMem[1034];
              ip = 1836;
        end

       1836 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1837;
              heapClock = ~ heapClock;
        end

       1837 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1035] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1838;
              heapClock = ~ heapClock;
        end

       1838 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[401] = localMem[1035];
              ip = 1839;
        end

       1839 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[401];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[400];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1840;
              heapClock = ~ heapClock;
        end

       1840 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1036] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1841;
              heapClock = ~ heapClock;
        end

       1841 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[402] = localMem[1036];
              ip = 1842;
        end

       1842 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[402] != localMem[362] ? 1883 : 1843;
        end

       1843 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1844;
              heapClock = ~ heapClock;
        end

       1844 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1037] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1845;
              heapClock = ~ heapClock;
        end

       1845 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[403] = localMem[1037];
              ip = 1846;
        end

       1846 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[403];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[375];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1847;
              heapClock = ~ heapClock;
        end

       1847 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1038] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1848;
              heapClock = ~ heapClock;
        end

       1848 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[404] = localMem[1038];
              ip = 1849;
        end

       1849 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1850;
              heapClock = ~ heapClock;
        end

       1850 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1039] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1851;
              heapClock = ~ heapClock;
        end

       1851 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[405] = localMem[1039];
              ip = 1852;
        end

       1852 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1040] = localMem[404];
              ip = 1853;
        end

       1853 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[405];                                                // Array to write to
              heapIndex   = localMem[400];                                                // Index of element to write to
              heapIn      = localMem[1040];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1854;
              heapClock = ~ heapClock;
        end

       1854 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1855;
              heapClock = ~ heapClock;
        end

       1855 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1041] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1856;
              heapClock = ~ heapClock;
        end

       1856 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[406] = localMem[1041];
              ip = 1857;
        end

       1857 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[406];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[375];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1858;
              heapClock = ~ heapClock;
        end

       1858 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1042] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1859;
              heapClock = ~ heapClock;
        end

       1859 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[407] = localMem[1042];
              ip = 1860;
        end

       1860 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1861;
              heapClock = ~ heapClock;
        end

       1861 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1043] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1862;
              heapClock = ~ heapClock;
        end

       1862 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[408] = localMem[1043];
              ip = 1863;
        end

       1863 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1044] = localMem[407];
              ip = 1864;
        end

       1864 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[408];                                                // Array to write to
              heapIndex   = localMem[400];                                                // Index of element to write to
              heapIn      = localMem[1044];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1865;
              heapClock = ~ heapClock;
        end

       1865 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1866;
              heapClock = ~ heapClock;
        end

       1866 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1045] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1867;
              heapClock = ~ heapClock;
        end

       1867 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[409] = localMem[1045];
              ip = 1868;
        end

       1868 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[375];
              heapArray  = localMem[409];
              ip = 1869;
              heapClock = ~ heapClock;
        end

       1869 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1870;
              heapClock = ~ heapClock;
        end

       1870 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1046] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1871;
              heapClock = ~ heapClock;
        end

       1871 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[410] = localMem[1046];
              ip = 1872;
        end

       1872 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[375];
              heapArray  = localMem[410];
              ip = 1873;
              heapClock = ~ heapClock;
        end

       1873 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[411] = localMem[400] + 1;
              ip = 1874;
        end

       1874 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1047] = localMem[411];
              ip = 1875;
        end

       1875 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[377];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1047];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1876;
              heapClock = ~ heapClock;
        end

       1876 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1877;
              heapClock = ~ heapClock;
        end

       1877 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1048] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1878;
              heapClock = ~ heapClock;
        end

       1878 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[412] = localMem[1048];
              ip = 1879;
        end

       1879 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1049] = localMem[378];
              ip = 1880;
        end

       1880 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[412];                                                // Array to write to
              heapIndex   = localMem[411];                                                // Index of element to write to
              heapIn      = localMem[1049];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1881;
              heapClock = ~ heapClock;
        end

       1881 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2176;
        end

       1882 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1882");
        end

       1883 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1883");
        end

       1884 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  1884");
        end

       1885 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1885");
        end

       1886 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1886");
        end

       1887 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1887");
        end

       1888 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1888");
        end

       1889 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1889");
        end

       1890 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1890");
        end

       1891 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1891");
        end

       1892 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1892");
        end

       1893 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1893");
        end

       1894 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1894");
        end

       1895 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1895");
        end

       1896 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1896");
        end

       1897 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1897");
        end

       1898 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1898");
        end

       1899 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1899");
        end

       1900 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1900");
        end

       1901 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1901");
        end

       1902 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1902");
        end

       1903 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1903");
        end

       1904 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1904");
        end

       1905 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1905");
        end

       1906 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1906");
        end

       1907 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1907");
        end

       1908 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1908");
        end

       1909 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1909");
        end

       1910 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1910");
        end

       1911 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1911");
        end

       1912 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1912");
        end

       1913 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1913");
        end

       1914 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1914");
        end

       1915 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1915");
        end

       1916 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1916");
        end

       1917 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1917");
        end

       1918 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1918");
        end

       1919 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1919");
        end

       1920 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1920");
        end

       1921 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1921");
        end

       1922 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1922");
        end

       1923 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1923");
        end

       1924 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1924");
        end

       1925 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1925");
        end

       1926 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1926");
        end

       1927 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1927");
        end

       1928 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1928");
        end

       1929 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1929");
        end

       1930 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1930");
        end

       1931 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1931");
        end

       1932 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1932");
        end

       1933 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1933");
        end

       1934 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1934");
        end

       1935 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1935");
        end

       1936 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1936");
        end

       1937 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1937");
        end

       1938 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1938");
        end

       1939 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1939");
        end

       1940 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1940");
        end

       1941 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1941");
        end

       1942 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1942");
        end

       1943 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1943");
        end

       1944 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1944");
        end

       1945 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1945");
        end

       1946 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1946");
        end

       1947 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1947");
        end

       1948 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1948");
        end

       1949 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1949");
        end

       1950 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1950");
        end

       1951 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1951");
        end

       1952 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1952");
        end

       1953 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1953");
        end

       1954 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1954");
        end

       1955 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1955");
        end

       1956 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1956");
        end

       1957 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1957");
        end

       1958 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1958");
        end

       1959 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1959");
        end

       1960 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1960");
        end

       1961 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1961");
        end

       1962 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1962");
        end

       1963 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1963");
        end

       1964 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1964");
        end

       1965 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1965");
        end

       1966 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1966");
        end

       1967 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1967");
        end

       1968 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1968");
        end

       1969 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1969");
        end

       1970 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1970");
        end

       1971 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1971");
        end

       1972 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1972");
        end

       1973 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1973");
        end

       1974 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1974");
        end

       1975 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1975");
        end

       1976 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1976");
        end

       1977 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1977");
        end

       1978 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1978");
        end

       1979 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1979");
        end

       1980 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1980");
        end

       1981 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1981");
        end

       1982 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1982");
        end

       1983 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1983");
        end

       1984 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1984");
        end

       1985 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1985");
        end

       1986 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1986");
        end

       1987 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1987");
        end

       1988 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1988");
        end

       1989 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1989");
        end

       1990 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1990");
        end

       1991 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1991");
        end

       1992 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1992");
        end

       1993 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1993");
        end

       1994 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1994");
        end

       1995 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1995");
        end

       1996 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1996");
        end

       1997 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1997");
        end

       1998 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1998");
        end

       1999 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1999");
        end

       2000 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2000");
        end

       2001 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2001");
        end

       2002 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2002");
        end

       2003 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2003");
        end

       2004 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2004");
        end

       2005 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2005");
        end

       2006 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2006");
        end

       2007 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2007");
        end

       2008 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2008");
        end

       2009 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2009");
        end

       2010 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2010");
        end

       2011 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2011");
        end

       2012 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2012");
        end

       2013 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2013");
        end

       2014 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2014");
        end

       2015 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2015");
        end

       2016 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2016");
        end

       2017 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2017");
        end

       2018 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2018");
        end

       2019 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2019");
        end

       2020 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2020");
        end

       2021 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2021");
        end

       2022 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2022");
        end

       2023 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2023");
        end

       2024 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2024");
        end

       2025 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2025");
        end

       2026 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2026");
        end

       2027 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2027");
        end

       2028 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2028");
        end

       2029 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2029");
        end

       2030 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2030");
        end

       2031 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2031");
        end

       2032 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2032");
        end

       2033 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2033");
        end

       2034 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2034");
        end

       2035 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2035");
        end

       2036 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2036");
        end

       2037 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2037");
        end

       2038 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2038");
        end

       2039 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2039");
        end

       2040 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2040");
        end

       2041 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2041");
        end

       2042 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2042");
        end

       2043 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2043");
        end

       2044 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2044");
        end

       2045 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2045");
        end

       2046 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2046");
        end

       2047 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2047");
        end

       2048 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2048");
        end

       2049 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2049");
        end

       2050 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2050");
        end

       2051 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2051");
        end

       2052 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2052");
        end

       2053 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2053");
        end

       2054 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2054");
        end

       2055 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2055");
        end

       2056 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2056");
        end

       2057 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2057");
        end

       2058 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2058");
        end

       2059 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2059");
        end

       2060 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2060");
        end

       2061 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2061");
        end

       2062 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2062");
        end

       2063 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2063");
        end

       2064 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2064");
        end

       2065 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2065");
        end

       2066 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2066");
        end

       2067 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2067");
        end

       2068 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2068");
        end

       2069 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2069");
        end

       2070 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2070");
        end

       2071 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2071");
        end

       2072 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2072");
        end

       2073 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2073");
        end

       2074 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2074");
        end

       2075 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2075");
        end

       2076 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2076");
        end

       2077 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2077");
        end

       2078 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2078");
        end

       2079 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2079");
        end

       2080 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2080");
        end

       2081 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2081");
        end

       2082 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2082");
        end

       2083 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2083");
        end

       2084 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2084");
        end

       2085 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2085");
        end

       2086 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2086");
        end

       2087 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2087");
        end

       2088 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2088");
        end

       2089 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2089");
        end

       2090 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2090");
        end

       2091 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2091");
        end

       2092 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2092");
        end

       2093 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2093");
        end

       2094 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2094");
        end

       2095 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2095");
        end

       2096 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2096");
        end

       2097 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2097");
        end

       2098 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2098");
        end

       2099 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2099");
        end

       2100 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2100");
        end

       2101 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2101");
        end

       2102 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2102");
        end

       2103 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2103");
        end

       2104 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2104");
        end

       2105 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2105");
        end

       2106 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2106");
        end

       2107 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2107");
        end

       2108 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2108");
        end

       2109 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2109");
        end

       2110 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2110");
        end

       2111 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2111");
        end

       2112 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2112");
        end

       2113 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2113");
        end

       2114 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2114");
        end

       2115 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2115");
        end

       2116 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2116");
        end

       2117 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2117");
        end

       2118 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2118");
        end

       2119 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2119");
        end

       2120 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2120");
        end

       2121 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2121");
        end

       2122 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2122");
        end

       2123 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2123");
        end

       2124 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2124");
        end

       2125 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2125");
        end

       2126 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2126");
        end

       2127 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2127");
        end

       2128 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2128");
        end

       2129 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2129");
        end

       2130 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2130");
        end

       2131 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2131");
        end

       2132 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2132");
        end

       2133 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2133");
        end

       2134 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2134");
        end

       2135 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2135");
        end

       2136 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2136");
        end

       2137 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2137");
        end

       2138 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2138");
        end

       2139 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2139");
        end

       2140 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2140");
        end

       2141 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2141");
        end

       2142 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2142");
        end

       2143 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2143");
        end

       2144 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2144");
        end

       2145 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2145");
        end

       2146 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2146");
        end

       2147 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2147");
        end

       2148 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2148");
        end

       2149 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2149");
        end

       2150 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2150");
        end

       2151 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2151");
        end

       2152 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2152");
        end

       2153 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2153");
        end

       2154 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2154");
        end

       2155 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2155");
        end

       2156 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2156");
        end

       2157 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2157");
        end

       2158 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2158");
        end

       2159 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2159");
        end

       2160 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2160");
        end

       2161 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2161");
        end

       2162 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2162");
        end

       2163 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2163");
        end

       2164 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2164");
        end

       2165 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2165");
        end

       2166 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2166");
        end

       2167 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2167");
        end

       2168 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2168");
        end

       2169 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2169");
        end

       2170 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2170");
        end

       2171 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2171");
        end

       2172 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2172");
        end

       2173 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2173");
        end

       2174 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2174");
        end

       2175 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2175");
        end

       2176 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2177;
        end

       2177 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[371] = 1;
              ip = 2178;
        end

       2178 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2181;
        end

       2179 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2180;
        end

       2180 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[371] = 0;
              ip = 2181;
        end

       2181 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2182;
        end

       2182 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2183;
        end

       2183 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2184;
        end

       2184 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2185;
        end

       2185 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[3];
              ip = 2186;
              heapClock = ~ heapClock;
        end

       2186 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2187;
        end

       2187 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1] = localMem[1] + 1;
              ip = 2188;
        end

       2188 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 14;
        end

       2189 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2190;
        end

       2190 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2191;
        end

       2191 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[478] = 0;
              ip = 2192;
        end

       2192 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2193;
        end

       2193 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[478] >= 66 ? 2301 : 2194;
        end

       2194 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[479] = localMem[478] + localMem[478];
              ip = 2195;
        end

       2195 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2196;
              heapClock = ~ heapClock;
        end

       2196 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[480] = heapOut;
              ip = 2197;
        end

       2197 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2198;
        end

       2198 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2199;
              heapClock = ~ heapClock;
        end

       2199 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1132] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2200;
              heapClock = ~ heapClock;
        end

       2200 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = localMem[1132];
              ip = 2201;
        end

       2201 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[481] != 0 ? 2209 : 2202;
        end

       2202 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2202");
        end

       2203 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2203");
        end

       2204 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2204");
        end

       2205 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2205");
        end

       2206 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2206");
        end

       2207 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2207");
        end

       2208 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2208");
        end

       2209 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2210;
        end

       2210 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2211;
        end

       2211 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[482] = 0;
              ip = 2212;
        end

       2212 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2213;
        end

       2213 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[482] >= 99 ? 2280 : 2214;
        end

       2214 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2215;
              heapClock = ~ heapClock;
        end

       2215 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1136] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2216;
              heapClock = ~ heapClock;
        end

       2216 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[483] = localMem[1136] - 1;
              ip = 2217;
        end

       2217 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2218;
              heapClock = ~ heapClock;
        end

       2218 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1137] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2219;
              heapClock = ~ heapClock;
        end

       2219 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[484] = localMem[1137];
              ip = 2220;
        end

       2220 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[484];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[483];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2221;
              heapClock = ~ heapClock;
        end

       2221 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1138] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2222;
              heapClock = ~ heapClock;
        end

       2222 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[478] <= localMem[1138] ? 2244 : 2223;
        end

       2223 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[485] = localMem[483] + 1;
              ip = 2224;
        end

       2224 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2225;
              heapClock = ~ heapClock;
        end

       2225 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1139] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2226;
              heapClock = ~ heapClock;
        end

       2226 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[486] = !localMem[1139];
              ip = 2227;
        end

       2227 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[486] == 0 ? 2235 : 2228;
        end

       2228 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2228");
        end

       2229 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2229");
        end

       2230 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2230");
        end

       2231 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2231");
        end

       2232 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2232");
        end

       2233 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2233");
        end

       2234 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2234");
        end

       2235 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2236;
        end

       2236 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2237;
              heapClock = ~ heapClock;
        end

       2237 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1143] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2238;
              heapClock = ~ heapClock;
        end

       2238 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[487] = localMem[1143];
              ip = 2239;
        end

       2239 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[487];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[485];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2240;
              heapClock = ~ heapClock;
        end

       2240 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1144] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2241;
              heapClock = ~ heapClock;
        end

       2241 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[488] = localMem[1144];
              ip = 2242;
        end

       2242 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = localMem[488];
              ip = 2243;
        end

       2243 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2277;
        end

       2244 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2245;
        end

       2245 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[478];
              heapAction = `Index;
              heapArray  = localMem[484];
              ip = 2246;
              heapClock = ~ heapClock;
        end

       2246 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[489] = heapOut;
              ip = 2247;
        end

       2247 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[489] == 0 ? 2255 : 2248;
        end

       2248 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1145] = localMem[481];
              ip = 2249;
        end

       2249 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[480];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1145];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2250;
              heapClock = ~ heapClock;
        end

       2250 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1146] = 1;
              ip = 2251;
        end

       2251 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[480];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1146];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2252;
              heapClock = ~ heapClock;
        end

       2252 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[1147] = localMem[489] - 1;
              ip = 2253;
        end

       2253 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[480];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1147];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2254;
              heapClock = ~ heapClock;
        end

       2254 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2284;
        end

       2255 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2256;
        end

       2256 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
              heapIn     = localMem[478];
              heapAction = `Less;
              heapArray  = localMem[484];
              ip = 2257;
              heapClock = ~ heapClock;
        end

       2257 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[490] = heapOut;
              ip = 2258;
        end

       2258 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2259;
              heapClock = ~ heapClock;
        end

       2259 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1148] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2260;
              heapClock = ~ heapClock;
        end

       2260 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[491] = !localMem[1148];
              ip = 2261;
        end

       2261 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[491] == 0 ? 2269 : 2262;
        end

       2262 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2262");
        end

       2263 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2263");
        end

       2264 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2264");
        end

       2265 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2265");
        end

       2266 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2266");
        end

       2267 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2267");
        end

       2268 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2268");
        end

       2269 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2270;
        end

       2270 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2271;
              heapClock = ~ heapClock;
        end

       2271 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1152] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2272;
              heapClock = ~ heapClock;
        end

       2272 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[492] = localMem[1152];
              ip = 2273;
        end

       2273 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[492];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[490];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2274;
              heapClock = ~ heapClock;
        end

       2274 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1153] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2275;
              heapClock = ~ heapClock;
        end

       2275 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[493] = localMem[1153];
              ip = 2276;
        end

       2276 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = localMem[493];
              ip = 2277;
        end

       2277 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2278;
        end

       2278 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[482] = localMem[482] + 1;
              ip = 2279;
        end

       2279 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2212;
        end

       2280 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2280");
        end

       2281 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  2281");
        end

       2282 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2282");
        end

       2283 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2283");
        end

       2284 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2285;
        end

       2285 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2286;
              heapClock = ~ heapClock;
        end

       2286 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1154] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2287;
              heapClock = ~ heapClock;
        end

       2287 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[494] = localMem[1154];
              ip = 2288;
        end

       2288 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2289;
              heapClock = ~ heapClock;
        end

       2289 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1155] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2290;
              heapClock = ~ heapClock;
        end

       2290 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[495] = localMem[1155];
              ip = 2291;
        end

       2291 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[494];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2292;
              heapClock = ~ heapClock;
        end

       2292 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1156] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2293;
              heapClock = ~ heapClock;
        end

       2293 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[496] = localMem[1156];
              ip = 2294;
        end

       2294 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[496];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[495];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2295;
              heapClock = ~ heapClock;
        end

       2295 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1157] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2296;
              heapClock = ~ heapClock;
        end

       2296 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[497] = localMem[1157];
              ip = 2297;
        end

       2297 :
        begin                                                                   // assertEq
          //$display("AAAA %4d %4d assertEq", steps, ip);
            ip = 2298;
        end

       2298 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2299;
        end

       2299 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[478] = localMem[478] + 1;
              ip = 2300;
        end

       2300 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2192;
        end

       2301 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2302;
        end

       2302 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2303;
              heapClock = ~ heapClock;
        end

       2303 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[498] = heapOut;
              ip = 2304;
        end

       2304 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2305;
        end

       2305 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2306;
              heapClock = ~ heapClock;
        end

       2306 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1158] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2307;
              heapClock = ~ heapClock;
        end

       2307 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[499] = localMem[1158];
              ip = 2308;
        end

       2308 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[499] != 0 ? 2316 : 2309;
        end

       2309 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2309");
        end

       2310 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2310");
        end

       2311 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2311");
        end

       2312 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2312");
        end

       2313 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2313");
        end

       2314 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2314");
        end

       2315 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2315");
        end

       2316 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2317;
        end

       2317 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2318;
        end

       2318 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[500] = 0;
              ip = 2319;
        end

       2319 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2320;
        end

       2320 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[500] >= 99 ? 2387 : 2321;
        end

       2321 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2322;
              heapClock = ~ heapClock;
        end

       2322 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1162] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2323;
              heapClock = ~ heapClock;
        end

       2323 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[501] = localMem[1162] - 1;
              ip = 2324;
        end

       2324 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2325;
              heapClock = ~ heapClock;
        end

       2325 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1163] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2326;
              heapClock = ~ heapClock;
        end

       2326 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[502] = localMem[1163];
              ip = 2327;
        end

       2327 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[502];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[501];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2328;
              heapClock = ~ heapClock;
        end

       2328 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1164] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2329;
              heapClock = ~ heapClock;
        end

       2329 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = -1 <= localMem[1164] ? 2351 : 2330;
        end

       2330 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2330");
        end

       2331 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2331");
        end

       2332 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2332");
        end

       2333 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  2333");
        end

       2334 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  2334");
        end

       2335 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2335");
        end

       2336 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2336");
        end

       2337 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2337");
        end

       2338 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2338");
        end

       2339 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2339");
        end

       2340 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2340");
        end

       2341 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2341");
        end

       2342 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2342");
        end

       2343 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2343");
        end

       2344 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2344");
        end

       2345 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2345");
        end

       2346 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2346");
        end

       2347 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2347");
        end

       2348 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2348");
        end

       2349 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2349");
        end

       2350 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2350");
        end

       2351 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2352;
        end

       2352 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = -1;
              heapAction = `Index;
              heapArray  = localMem[502];
              ip = 2353;
              heapClock = ~ heapClock;
        end

       2353 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[507] = heapOut;
              ip = 2354;
        end

       2354 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[507] == 0 ? 2362 : 2355;
        end

       2355 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2355");
        end

       2356 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2356");
        end

       2357 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2357");
        end

       2358 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2358");
        end

       2359 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  2359");
        end

       2360 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2360");
        end

       2361 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2361");
        end

       2362 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2363;
        end

       2363 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
              heapIn     = -1;
              heapAction = `Less;
              heapArray  = localMem[502];
              ip = 2364;
              heapClock = ~ heapClock;
        end

       2364 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[508] = heapOut;
              ip = 2365;
        end

       2365 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2366;
              heapClock = ~ heapClock;
        end

       2366 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1174] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2367;
              heapClock = ~ heapClock;
        end

       2367 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[509] = !localMem[1174];
              ip = 2368;
        end

       2368 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[509] == 0 ? 2376 : 2369;
        end

       2369 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1175] = localMem[499];
              ip = 2370;
        end

       2370 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[498];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1175];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2371;
              heapClock = ~ heapClock;
        end

       2371 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1176] = 0;
              ip = 2372;
        end

       2372 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[498];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1176];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2373;
              heapClock = ~ heapClock;
        end

       2373 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1177] = localMem[508];
              ip = 2374;
        end

       2374 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[498];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1177];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2375;
              heapClock = ~ heapClock;
        end

       2375 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2391;
        end

       2376 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2377;
        end

       2377 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2378;
              heapClock = ~ heapClock;
        end

       2378 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1178] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2379;
              heapClock = ~ heapClock;
        end

       2379 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[510] = localMem[1178];
              ip = 2380;
        end

       2380 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[510];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[508];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2381;
              heapClock = ~ heapClock;
        end

       2381 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1179] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2382;
              heapClock = ~ heapClock;
        end

       2382 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[511] = localMem[1179];
              ip = 2383;
        end

       2383 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[499] = localMem[511];
              ip = 2384;
        end

       2384 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2385;
        end

       2385 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[500] = localMem[500] + 1;
              ip = 2386;
        end

       2386 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2319;
        end

       2387 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2387");
        end

       2388 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  2388");
        end

       2389 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2389");
        end

       2390 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2390");
        end

       2391 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2392;
        end

       2392 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2393;
              heapClock = ~ heapClock;
        end

       2393 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1180] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2394;
              heapClock = ~ heapClock;
        end

       2394 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[512] = localMem[1180];
              ip = 2395;
        end

       2395 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
            ip = 2396;
        end

       2396 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2397;
              heapClock = ~ heapClock;
        end

       2397 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[513] = heapOut;
              ip = 2398;
        end

       2398 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2399;
        end

       2399 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2400;
              heapClock = ~ heapClock;
        end

       2400 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1181] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2401;
              heapClock = ~ heapClock;
        end

       2401 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[514] = localMem[1181];
              ip = 2402;
        end

       2402 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[514] != 0 ? 2410 : 2403;
        end

       2403 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2403");
        end

       2404 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2404");
        end

       2405 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2405");
        end

       2406 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2406");
        end

       2407 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2407");
        end

       2408 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2408");
        end

       2409 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2409");
        end

       2410 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2411;
        end

       2411 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2412;
        end

       2412 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[515] = 0;
              ip = 2413;
        end

       2413 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2414;
        end

       2414 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[515] >= 99 ? 2481 : 2415;
        end

       2415 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[514];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2416;
              heapClock = ~ heapClock;
        end

       2416 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1185] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2417;
              heapClock = ~ heapClock;
        end

       2417 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[516] = localMem[1185] - 1;
              ip = 2418;
        end

       2418 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[514];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2419;
              heapClock = ~ heapClock;
        end

       2419 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1186] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2420;
              heapClock = ~ heapClock;
        end

       2420 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[517] = localMem[1186];
              ip = 2421;
        end

       2421 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[517];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[516];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2422;
              heapClock = ~ heapClock;
        end

       2422 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1187] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2423;
              heapClock = ~ heapClock;
        end

       2423 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = 66 <= localMem[1187] ? 2445 : 2424;
        end

       2424 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[518] = localMem[516] + 1;
              ip = 2425;
        end

       2425 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[514];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2426;
              heapClock = ~ heapClock;
        end

       2426 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1188] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2427;
              heapClock = ~ heapClock;
        end

       2427 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[519] = !localMem[1188];
              ip = 2428;
        end

       2428 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[519] == 0 ? 2436 : 2429;
        end

       2429 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1189] = localMem[514];
              ip = 2430;
        end

       2430 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[513];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1189];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2431;
              heapClock = ~ heapClock;
        end

       2431 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1190] = 2;
              ip = 2432;
        end

       2432 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[513];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1190];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2433;
              heapClock = ~ heapClock;
        end

       2433 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1191] = localMem[518];
              ip = 2434;
        end

       2434 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[513];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1191];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2435;
              heapClock = ~ heapClock;
        end

       2435 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2485;
        end

       2436 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2437;
        end

       2437 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[514];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2438;
              heapClock = ~ heapClock;
        end

       2438 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1192] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2439;
              heapClock = ~ heapClock;
        end

       2439 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[520] = localMem[1192];
              ip = 2440;
        end

       2440 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[520];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[518];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2441;
              heapClock = ~ heapClock;
        end

       2441 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1193] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2442;
              heapClock = ~ heapClock;
        end

       2442 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[521] = localMem[1193];
              ip = 2443;
        end

       2443 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[514] = localMem[521];
              ip = 2444;
        end

       2444 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2478;
        end

       2445 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2445");
        end

       2446 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  2446");
        end

       2447 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2447");
        end

       2448 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  2448");
        end

       2449 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2449");
        end

       2450 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2450");
        end

       2451 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2451");
        end

       2452 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2452");
        end

       2453 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  2453");
        end

       2454 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2454");
        end

       2455 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2455");
        end

       2456 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2456");
        end

       2457 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed  2457");
        end

       2458 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2458");
        end

       2459 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2459");
        end

       2460 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2460");
        end

       2461 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  2461");
        end

       2462 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  2462");
        end

       2463 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2463");
        end

       2464 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2464");
        end

       2465 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2465");
        end

       2466 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2466");
        end

       2467 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2467");
        end

       2468 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2468");
        end

       2469 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2469");
        end

       2470 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2470");
        end

       2471 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2471");
        end

       2472 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2472");
        end

       2473 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2473");
        end

       2474 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2474");
        end

       2475 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2475");
        end

       2476 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2476");
        end

       2477 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2477");
        end

       2478 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2479;
        end

       2479 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[515] = localMem[515] + 1;
              ip = 2480;
        end

       2480 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2413;
        end

       2481 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2481");
        end

       2482 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  2482");
        end

       2483 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2483");
        end

       2484 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2484");
        end

       2485 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2486;
        end

       2486 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[513];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2487;
              heapClock = ~ heapClock;
        end

       2487 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1203] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2488;
              heapClock = ~ heapClock;
        end

       2488 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[527] = localMem[1203];
              ip = 2489;
        end

       2489 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
            ip = 2490;
        end
      endcase
      success  = 1;
      finished = steps >  36159;
    end
  end

endmodule
