// Check double frees, over allocation
// Check access to unallocated arrays or elements
// Check push overflow, pop underflow
// Next Message 10000280
`define Reset        1  /* Zero all memory sizes                               */
`define Write        2  /* Write an element                                    */
`define Read         3  /* Read an element                                     */
`define Size         4  /* Size of array                                       */
`define Inc          5  /* Increment size of array if possible                 */
`define Dec          6  /* Decrement size of array if possible                 */
`define Index        7  /* Index of element in array                           */
`define Less         8  /* Elements of array less than in                      */
`define Greater      9  /* Elements of array greater than in                   */
`define Up          10  /* Move array up                                       */
`define Down        11  /* Move array down                                     */
`define Long1       12  /* Move long first step                                */
`define Long2       13  /* Move long last  step                                */
`define Push        14  /* Push if possible                                    */
`define Pop         15  /* Pop if possible                                     */
`define Dump        16  /* Dump                                                */
`define Resize      17  /* Resize an array                                     */
`define Alloc       18  /* Allocate a new array before using it                */
`define Free        19  /* Free an array for reuse                             */
`define Add         20  /* Add to an element returning the new value           */
`define AddAfter    21  /* Add to an element returning the previous value      */
`define Subtract    22  /* Subtract to an element returning the new value      */
`define SubAfter    23  /* Subtract to an element returning the previous value */
`define ShiftLeft   24  /* Shift left                                          */
`define ShiftRight  25  /* Shift right                                         */
`define NotLogical  26  /* Not - logical                                       */
`define Not         27  /* Not - bitwise                                       */
`define Or          28  /* Or                                                  */
`define Xor         29  /* Xor                                                 */
`define And         30  /* And                                                 */

module Memory
#(parameter integer ADDRESS_BITS =  8,                                          // Number of bits in an address
  parameter integer INDEX_BITS   =  3,                                          // Bits in in an index
  parameter integer DATA_BITS    = 16)                                          // Width of an element in bits
 (input wire                    clock,                                          // Clock to drive array operations
  input wire[7:0]               action,                                         // Operation to be performed on array
  input wire [ADDRESS_BITS-1:0] array,                                          // The number of the array to work on
  input wire [INDEX_BITS  -1:0] index,                                          // Index within array
  input wire [DATA_BITS   -1:0] in,                                             // Input data
  output reg [DATA_BITS   -1:0] out,                                            // Output data
  output reg [31:0]             error);                                         // Error

  parameter integer ARRAY_LENGTH = 2**INDEX_BITS;                               // Maximum index
  parameter integer ARRAYS       = 2**ADDRESS_BITS;                             // Number of memory elements for both arrays and elements

  reg [DATA_BITS   -1:0] memory     [ARRAYS-1:0][ARRAY_LENGTH-1:0];             // Memory containing arrays in fixed blocks
  reg [DATA_BITS   -1:0] copy                   [ARRAY_LENGTH-1:0];             // Copy of one array
  reg [INDEX_BITS    :0] arraySizes [ARRAYS-1:0];                               // Current size of each array
  reg [ADDRESS_BITS-1:0] freedArrays[ARRAYS-1:0];                               // Currently freed arrays
  reg                    allocations[ARRAYS-1:0];                               // Currently allocated arrays

  integer allocatedArrays;                                                      // Arrays allocated
  integer freedArraysTop;                                                       // Top of the freed arrays stack
  integer result;                                                               // Result of each array operation
  integer size;                                                                 // Size of current array
  integer moveLongStartArray;                                                   // Source array of move long
  integer moveLongStartIndex;                                                   // Source index of move long
  integer i, a, b;                                                              // Index

  task checkWriteable(input integer err);                                       // Check a memory is writable
    begin
       error = 0;
       if (array >= allocatedArrays) begin
         //$display("Array has not been allocated, array %d", array);
         error = err;
       end
       if (!allocations[array]) begin
         //$display("Array has been freed, array %d", array);
         error = err + 1;
       end
    end
  endtask

  task checkReadable(input integer err);                                        // Check a memory locationis readable
    begin
       checkWriteable(err);
       if (index >= arraySizes[array]) begin
         //$display("Access outside array bounds, array %d, size: %d, access: %d", array, arraySizes[array], index);
         error = err + 2;
       end
    end
  endtask

  task dump;                                                                    // Dump some memory
    begin
      //$display("    %2d %2d %2d", arraySizes[0], arraySizes[1], arraySizes[2]);
      for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
        //$display("%2d  %2d %2d %2d", i, memory[0][i], memory[1][i], memory[2][i]);
      end
      //$display("    %2d %2d %2d", allocations[0], allocations[1], allocations[2]);
    end
  endtask

  always @(posedge clock) begin                                                 // Each transition
    case(action)                                                                // Decode request
      `Reset: begin                                                             // Reset
        freedArraysTop = 0;                                                     // Free all arrays
        allocatedArrays = 0;
      end

      `Write: begin                                                             // Write
        checkWriteable(10000010);
        if (!error) begin
          memory[array][index] = in;
          if (index >= arraySizes[array] && index < ARRAY_LENGTH) begin
            arraySizes[array] = index + 1;
          end
          out = in;
        end
      end

      `Read: begin                                                              // Read
        checkReadable(10000020);
        if (!error) begin
          out = memory[array][index];
        end
      end

      `Size: begin                                                              // Size
        checkWriteable(10000030);
        if (!error) begin
          out = arraySizes[array];
        end
      end

      `Dec: begin                                                               // Decrement
        checkWriteable(10000040);
        if (!error) begin
          if (arraySizes[array] > 0) arraySizes[array] = arraySizes[array] - 1;
          else begin
            //$display("Attempt to decrement empty array, array %d", array); error = 10000044;
          end
        end
      end

      `Inc: begin                                                               // Increment
        checkWriteable(10000050);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;
          else begin
            //$display("Attempt to decrement full array, array %d", array);  error = 10000054;
          end
        end
      end

      `Index: begin                                                             // Index
        checkWriteable(10000060);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] == in) result = i + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Less: begin                                                              // Count less
        checkWriteable(10000070);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] < in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Greater: begin                                                           // Count greater
        checkWriteable(10000080);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] > in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Down: begin                                                              // Down
        checkWriteable(10000270);
        if (!error) begin
          size   = arraySizes[array];
          if (size > 0) begin
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i]; // Copy source array
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                       // Move original array up
              if (i > index && i <= size) begin
                memory[array][i-1] = copy[i];
              end
            end
            out = copy[index];                                                  // Return replaced value
            arraySizes[array] = arraySizes[array] - 1;                          // Decrease array size
          end
          else error = 100000274;                                               // Orignal array was emoty so we cannot shift it down
        end
      end

      `Up: begin                                                                // Up
        checkWriteable(10000090);
        if (!error) begin
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i];   // Copy source array
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Move original array up
            if (i > index && i <= size) begin
              memory[array][i] = copy[i-1];
            end
          end
          memory[array][index] = in;                                            // Insert new value
          if (size < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;   // Increase array size
        end
      end

      `Long1: begin                                                             // Move long start
        checkReadable(10000100);
        if (!error) begin
          moveLongStartArray = array;                                           // Record source
          moveLongStartIndex = index;
        end
      end

      `Long2: begin                                                             // Move long finish
        checkWriteable(10000110);
        if (!error) begin
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Copy from source to target
            if (i < in && index + i < ARRAY_LENGTH && moveLongStartIndex+i < ARRAY_LENGTH) begin
              memory[array][index+i] = memory[moveLongStartArray][moveLongStartIndex+i];
              if (index+i >= arraySizes[array]) arraySizes[array] = index+i+1;
            end
          end
        end
      end

      `Push: begin                                                              // Push
        checkWriteable(10000120);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) begin
            memory[array][arraySizes[array]] = in;
            arraySizes[array] = arraySizes[array] + 1;
          end
          else begin
            //$display("Attempt to push to full array, array %d, value %d", array, in);  error = 10000124;
          end
        end
      end

      `Pop: begin                                                               // Pop
        checkWriteable(10000130);
        if (!error) begin
          if (arraySizes[array] > 0) begin
            arraySizes[array] = arraySizes[array] - 1;
            out = memory[array][arraySizes[array]];
          end
          else begin
            //$display("Attempt to pop empty array, array %d", array); error = 10000134;
          end
        end
      end

      `Dump: begin                                                              // Dump
        dump();
      end

      `Resize: begin                                                            // Resize
        checkWriteable(10000140);
        if (!error) begin
          if (in <= ARRAY_LENGTH) arraySizes[array] = in;
          else begin
            //$display("Attempt to make an array too large, array %d, max %d, size %d", array, ARRAY_LENGTH, in); error = 10000144;
          end
        end
      end

      `Alloc: begin                                                             // Allocate an array
        if (freedArraysTop > 0) begin                                           // Reuse a freed array
          freedArraysTop = freedArraysTop - 1;
          result = freedArrays[freedArraysTop];
        end
        else if (allocatedArrays < ARRAYS-1) begin                              // Allocate a new array - assumes enough memory
          result          = allocatedArrays;
          allocatedArrays = allocatedArrays + 1;
        end
        else begin
          //$display("Out of memory, cannot allocate a new array"); error = 10000270;
        end
        allocations[result] = 1;                                                // Allocated
        arraySizes[result] = 0;                                                 // Empty array
        out = result;
      end

      `Free: begin                                                              // Free an array
        checkWriteable(10000150);
        if (!error) begin
          freedArrays[freedArraysTop] = array;                                  // Relies on the user not re freeing a freed array - we should probably hve another array to prevent this
          allocations[array]          = 0;                                      // No longer allocated
          freedArraysTop = freedArraysTop + 1;
        end
      end

      `Add: begin                                                               // Add to an element
        checkReadable(10000160);
        if (!error) begin
          memory[array][index] = memory[array][index] + in;
          out = memory[array][index];
        end
      end

      `AddAfter: begin                                                          // Add to an element after putting the content of the element on out
        checkReadable(10000170);
        if (!error) begin
        out = memory[array][index];
        memory[array][index] = memory[array][index] + in;
        end
      end

      `Subtract: begin                                                          // Subtract from an element
        checkReadable(10000180);
        if (!error) begin
          memory[array][index] = memory[array][index] - in;
          out = memory[array][index];
        end
      end

      `SubAfter: begin                                                          // Subtract from an element after putting the content of the element on out
        checkReadable(10000190);
        if (!error) begin
          out = memory[array][index];
          memory[array][index] = memory[array][index] - in;
        end
      end

      `ShiftLeft: begin                                                         // Shift left
        checkReadable(10000200);
        if (!error) begin
          memory[array][index] = memory[array][index] << in;
          out = memory[array][index];
        end
      end

      `ShiftRight: begin                                                        // Shift right
        checkReadable(10000210);
        if (!error) begin
          memory[array][index] = memory[array][index] >> in;
          out = memory[array][index];
        end
      end

      `NotLogical: begin                                                        // Not logical
        checkReadable(10000220);
        if (!error) begin
          memory[array][index] = !memory[array][index];
          out = memory[array][index];
        end
      end

      `Not: begin                                                               // Not
        checkReadable(10000230);
        if (!error) begin
          memory[array][index] = ~memory[array][index];
          out = memory[array][index];
        end
      end

      `Or: begin                                                                // Or
        checkReadable(10000240);
        if (!error) begin
          memory[array][index] = memory[array][index] | in;
          out = memory[array][index];
        end
      end

      `Xor: begin                                                               // Xor
        checkReadable(10000250);
        if (!error) begin
          memory[array][index] = memory[array][index] ^ in;
          out = memory[array][index];
        end
      end

      `And: begin                                                               // And
        checkReadable(10000260);
        if (!error) begin
          memory[array][index] = memory[array][index] & in;
          out = memory[array][index];
        end
      end
    endcase
  end
endmodule
//-----------------------------------------------------------------------------
// Fpga test
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga                                                                     // Run test programs
 (input  wire clock,                                                            // Driving clock
  input  wire reset,                                                            // Restart program
  output reg  finished,                                                         // Goes high when the program has finished
  output reg  success);                                                         // Goes high on finish if all the tests passed

  reg                heapClock;                                                 // Clock to drive array operations
  reg [7:0]          heapAction;                                                // Operation to be performed on array
  reg [       9-1:0] heapArray;                                         // The number of the array to work on
  reg [       3-1:0] heapIndex;                                         // Index within array
  reg [      12-1:0] heapIn;                                            // Input data
  reg [      12-1:0] heapOut;                                           // Output data
  reg [31        :0] heapError;                                                 // Error on heap operation if not zero

  Memory                                                                        // Memory module
   #(       9,        3,       12)                          // Address bits, index bits, data bits
    heap(                                                                       // Create heap memory
    .clock  (heapClock),
    .action (heapAction),
    .array  (heapArray),
    .index  (heapIndex),
    .in     (heapIn),
    .out    (heapOut),
    .error  (heapError)
  );
  reg [      12-1:0] localMem[    1165-1:0];                       // Local memory
  reg [      12-1:0]   outMem[      67  -1:0];                       // Out channel
  reg [      12-1:0]    inMem[       1   -1:0];                       // In channel

  integer inMemPos;                                                             // Current position in input channel
  integer outMemPos;                                                            // Position in output channel

  integer ip;                                                                   // Instruction pointer
  integer steps;                                                                // Number of steps executed so far
  integer i, j, k;                                                              // A useful counter

  always @(posedge clock) begin                                                 // Each instruction
    if (reset) begin
      ip             = 0;
      steps          = 0;
      inMemPos       = 0;
      outMemPos      = 0;
      finished       = 0;
      success        = 0;

    end
    else begin
      case(ip)

          0 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1;
        end

          1 :
        begin                                                                   // start
          //$display("AAAA %4d %4d start", steps, ip);
              heapAction = `Reset;                                              // Reset heap memory
              ip = 2;
              heapClock = 1;
        end

          2 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3;
        end

          3 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 4;
              heapClock = 1;
        end

          4 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[0] = heapOut;
              ip = 5;
        end

          5 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 6;
        end

          6 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[512] = 3;
              ip = 7;
        end

          7 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[512];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 8;
              heapClock = 1;
        end

          8 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 9;
        end

          9 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[513] = 0;
              ip = 10;
        end

         10 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[513];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 11;
              heapClock = 1;
        end

         11 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 12;
        end

         12 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[514] = 0;
              ip = 13;
        end

         13 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[514];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 14;
              heapClock = 1;
        end

         14 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 15;
        end

         15 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[515] = 0;
              ip = 16;
        end

         16 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[515];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 17;
              heapClock = 1;
        end

         17 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 18;
        end

         18 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 19;
        end

         19 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1] = 0;
              ip = 20;
        end

         20 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 21;
        end

         21 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[1] >= 66 ? 3248 : 22;
        end

         22 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[2] = localMem[1] + localMem[1];
              ip = 23;
        end

         23 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 24;
              heapClock = 1;
        end

         24 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[3] = heapOut;
              ip = 25;
        end

         25 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 26;
        end

         26 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 27;
        end

         27 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 28;
              heapClock = 1;
        end

         28 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 29;
        end

         29 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[516] = heapOut;                                                     // Data retrieved from heap memory
              ip = 30;
              heapClock = 1;
        end

         30 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 31;
        end

         31 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[4] = localMem[516];
              ip = 32;
        end

         32 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[4] != 0 ? 113 : 33;
        end

         33 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 34;
              heapClock = 1;
        end

         34 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[5] = heapOut;
              ip = 35;
        end

         35 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 36;
        end

         36 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[517] = 1;
              ip = 37;
        end

         37 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[517];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 38;
              heapClock = 1;
        end

         38 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 39;
        end

         39 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[518] = 0;
              ip = 40;
        end

         40 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[518];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 41;
              heapClock = 1;
        end

         41 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 42;
        end

         42 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 43;
              heapClock = 1;
        end

         43 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[6] = heapOut;
              ip = 44;
        end

         44 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 45;
        end

         45 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[519] = localMem[6];
              ip = 46;
        end

         46 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[519];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 47;
              heapClock = 1;
        end

         47 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 48;
        end

         48 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 49;
              heapClock = 1;
        end

         49 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[7] = heapOut;
              ip = 50;
        end

         50 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 51;
        end

         51 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[520] = localMem[7];
              ip = 52;
        end

         52 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[520];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 53;
              heapClock = 1;
        end

         53 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 54;
        end

         54 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[521] = 0;
              ip = 55;
        end

         55 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[521];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 56;
              heapClock = 1;
        end

         56 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 57;
        end

         57 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[522] = localMem[0];
              ip = 58;
        end

         58 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[522];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 59;
              heapClock = 1;
        end

         59 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 60;
        end

         60 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 61;
              heapClock = 1;
        end

         61 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 62;
        end

         62 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[523] = heapOut;                                                     // Data retrieved from heap memory
              ip = 63;
              heapClock = 1;
        end

         63 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 64;
        end

         64 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[524] = localMem[523] + 1;
              ip = 65;
        end

         65 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[524];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 66;
              heapClock = 1;
        end

         66 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 67;
        end

         67 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 68;
              heapClock = 1;
        end

         68 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 69;
        end

         69 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[525] = heapOut;                                                     // Data retrieved from heap memory
              ip = 70;
              heapClock = 1;
        end

         70 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 71;
        end

         71 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[526] = localMem[525];
              ip = 72;
        end

         72 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[5];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[526];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 73;
              heapClock = 1;
        end

         73 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 74;
        end

         74 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 75;
              heapClock = 1;
        end

         75 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 76;
        end

         76 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[527] = heapOut;                                                     // Data retrieved from heap memory
              ip = 77;
              heapClock = 1;
        end

         77 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 78;
        end

         78 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[8] = localMem[527];
              ip = 79;
        end

         79 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[528] = localMem[1];
              ip = 80;
        end

         80 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[8];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[528];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 81;
              heapClock = 1;
        end

         81 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 82;
        end

         82 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 83;
              heapClock = 1;
        end

         83 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 84;
        end

         84 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[529] = heapOut;                                                     // Data retrieved from heap memory
              ip = 85;
              heapClock = 1;
        end

         85 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 86;
        end

         86 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[9] = localMem[529];
              ip = 87;
        end

         87 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[530] = localMem[2];
              ip = 88;
        end

         88 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[9];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[530];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 89;
              heapClock = 1;
        end

         89 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 90;
        end

         90 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 91;
              heapClock = 1;
        end

         91 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 92;
        end

         92 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[531] = heapOut;                                                     // Data retrieved from heap memory
              ip = 93;
              heapClock = 1;
        end

         93 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 94;
        end

         94 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[532] = localMem[531] + 1;
              ip = 95;
        end

         95 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[532];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 96;
              heapClock = 1;
        end

         96 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 97;
        end

         97 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[533] = localMem[5];
              ip = 98;
        end

         98 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[533];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 99;
              heapClock = 1;
        end

         99 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 100;
        end

        100 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 101;
              heapClock = 1;
        end

        101 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 102;
        end

        102 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[534] = heapOut;                                                     // Data retrieved from heap memory
              ip = 103;
              heapClock = 1;
        end

        103 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 104;
        end

        104 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[10] = localMem[534];
              ip = 105;
        end

        105 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[10];
              ip = 106;
              heapClock = 1;
        end

        106 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[5];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 107;
              heapClock = 1;
        end

        107 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 108;
        end

        108 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[535] = heapOut;                                                     // Data retrieved from heap memory
              ip = 109;
              heapClock = 1;
        end

        109 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 110;
        end

        110 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[11] = localMem[535];
              ip = 111;
        end

        111 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[11];
              ip = 112;
              heapClock = 1;
        end

        112 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3243;
        end

        113 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 114;
        end

        114 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 115;
              heapClock = 1;
        end

        115 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 116;
        end

        116 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[536] = heapOut;                                                     // Data retrieved from heap memory
              ip = 117;
              heapClock = 1;
        end

        117 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 118;
        end

        118 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[12] = localMem[536];
              ip = 119;
        end

        119 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 120;
              heapClock = 1;
        end

        120 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 121;
        end

        121 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[537] = heapOut;                                                     // Data retrieved from heap memory
              ip = 122;
              heapClock = 1;
        end

        122 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 123;
        end

        123 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[13] = localMem[537];
              ip = 124;
        end

        124 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[12] >= localMem[13] ? 228 : 125;
        end

        125 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 126;
              heapClock = 1;
        end

        126 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 127;
        end

        127 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[538] = heapOut;                                                     // Data retrieved from heap memory
              ip = 128;
              heapClock = 1;
        end

        128 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 129;
        end

        129 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[14] = localMem[538];
              ip = 130;
        end

        130 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[14] != 0 ? 227 : 131;
        end

        131 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 132;
              heapClock = 1;
        end

        132 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 133;
        end

        133 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[539] = heapOut;                                                     // Data retrieved from heap memory
              ip = 134;
              heapClock = 1;
        end

        134 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 135;
        end

        135 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[15] = !localMem[539];
              ip = 136;
        end

        136 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[15] == 0 ? 226 : 137;
        end

        137 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 138;
              heapClock = 1;
        end

        138 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 139;
        end

        139 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[540] = heapOut;                                                     // Data retrieved from heap memory
              ip = 140;
              heapClock = 1;
        end

        140 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 141;
        end

        141 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[16] = localMem[540];
              ip = 142;
        end

        142 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[1];
              heapAction = `Index;
              heapArray  = localMem[16];
              ip = 143;
              heapClock = 1;
        end

        143 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[17] = heapOut;
              ip = 144;
        end

        144 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 145;
        end

        145 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[17] == 0 ? 156 : 146;
        end

        146 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   146");
        end

        147 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   147");
        end

        148 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   148");
        end

        149 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   149");
        end

        150 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   150");
        end

        151 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   151");
        end

        152 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   152");
        end

        153 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   153");
        end

        154 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   154");
        end

        155 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   155");
        end

        156 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 157;
        end

        157 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[12];
              heapArray  = localMem[16];
              ip = 158;
              heapClock = 1;
        end

        158 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 159;
              heapClock = 1;
        end

        159 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 160;
        end

        160 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[543] = heapOut;                                                     // Data retrieved from heap memory
              ip = 161;
              heapClock = 1;
        end

        161 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 162;
        end

        162 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[19] = localMem[543];
              ip = 163;
        end

        163 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[12];
              heapArray  = localMem[19];
              ip = 164;
              heapClock = 1;
        end

        164 :
        begin                                                                   // arrayCountGreater
          //$display("AAAA %4d %4d arrayCountGreater", steps, ip);
              heapIn     = localMem[1];
              heapAction = `Greater;
              heapArray  = localMem[16];
              ip = 165;
              heapClock = 1;
        end

        165 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[20] = heapOut;
              ip = 166;
        end

        166 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 167;
        end

        167 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[20] != 0 ? 195 : 168;
        end

        168 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 169;
              heapClock = 1;
        end

        169 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 170;
        end

        170 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[544] = heapOut;                                                     // Data retrieved from heap memory
              ip = 171;
              heapClock = 1;
        end

        171 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 172;
        end

        172 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[21] = localMem[544];
              ip = 173;
        end

        173 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[545] = localMem[1];
              ip = 174;
        end

        174 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[21];                                                // Array to write to
              heapIndex   = localMem[12];                                                // Index of element to write to
              heapIn      = localMem[545];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 175;
              heapClock = 1;
        end

        175 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 176;
        end

        176 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[4];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 177;
              heapClock = 1;
        end

        177 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 178;
        end

        178 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[546] = heapOut;                                                     // Data retrieved from heap memory
              ip = 179;
              heapClock = 1;
        end

        179 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 180;
        end

        180 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[22] = localMem[546];
              ip = 181;
        end

        181 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[547] = localMem[2];
              ip = 182;
        end

        182 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[22];                                                // Array to write to
              heapIndex   = localMem[12];                                                // Index of element to write to
              heapIn      = localMem[547];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 183;
              heapClock = 1;
        end

        183 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 184;
        end

        184 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[548] = localMem[12] + 1;
              ip = 185;
        end

        185 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[4];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[548];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 186;
              heapClock = 1;
        end

        186 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 187;
        end

        187 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 188;
              heapClock = 1;
        end

        188 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 189;
        end

        189 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[549] = heapOut;                                                     // Data retrieved from heap memory
              ip = 190;
              heapClock = 1;
        end

        190 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 191;
        end

        191 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[550] = localMem[549] + 1;
              ip = 192;
        end

        192 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[550];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 193;
              heapClock = 1;
        end

        193 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 194;
        end

        194 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3243;
        end

        195 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   195");
        end

        196 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed   196");
        end

        197 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   197");
        end

        198 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   198");
        end

        199 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   199");
        end

        200 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   200");
        end

        201 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   201");
        end

        202 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   202");
        end

        203 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   203");
        end

        204 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   204");
        end

        205 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   205");
        end

        206 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   206");
        end

        207 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   207");
        end

        208 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   208");
        end

        209 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   209");
        end

        210 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   210");
        end

        211 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   211");
        end

        212 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   212");
        end

        213 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   213");
        end

        214 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   214");
        end

        215 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   215");
        end

        216 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   216");
        end

        217 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   217");
        end

        218 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   218");
        end

        219 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   219");
        end

        220 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   220");
        end

        221 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   221");
        end

        222 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   222");
        end

        223 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   223");
        end

        224 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   224");
        end

        225 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   225");
        end

        226 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 227;
        end

        227 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 228;
        end

        228 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 229;
        end

        229 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 230;
              heapClock = 1;
        end

        230 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 231;
        end

        231 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[557] = heapOut;                                                     // Data retrieved from heap memory
              ip = 232;
              heapClock = 1;
        end

        232 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 233;
        end

        233 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[26] = localMem[557];
              ip = 234;
        end

        234 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 235;
        end

        235 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 236;
              heapClock = 1;
        end

        236 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 237;
        end

        237 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[558] = heapOut;                                                     // Data retrieved from heap memory
              ip = 238;
              heapClock = 1;
        end

        238 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 239;
        end

        239 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[28] = localMem[558];
              ip = 240;
        end

        240 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 241;
              heapClock = 1;
        end

        241 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 242;
        end

        242 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[559] = heapOut;                                                     // Data retrieved from heap memory
              ip = 243;
              heapClock = 1;
        end

        243 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 244;
        end

        244 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[29] = localMem[559];
              ip = 245;
        end

        245 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 246;
              heapClock = 1;
        end

        246 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 247;
        end

        247 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[560] = heapOut;                                                     // Data retrieved from heap memory
              ip = 248;
              heapClock = 1;
        end

        248 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 249;
        end

        249 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[30] = localMem[560];
              ip = 250;
        end

        250 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[28] <  localMem[30] ? 935 : 251;
        end

        251 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[31] = localMem[30];
              ip = 252;
        end

        252 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[31] = localMem[31] >> 1;
              ip = 253;
              ip = 253;
        end

        253 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[32] = localMem[31] + 1;
              ip = 254;
        end

        254 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 255;
              heapClock = 1;
        end

        255 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 256;
        end

        256 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[561] = heapOut;                                                     // Data retrieved from heap memory
              ip = 257;
              heapClock = 1;
        end

        257 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 258;
        end

        258 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[33] = localMem[561];
              ip = 259;
        end

        259 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[33] == 0 ? 565 : 260;
        end

        260 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   260");
        end

        261 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   261");
        end

        262 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   262");
        end

        263 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   263");
        end

        264 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   264");
        end

        265 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   265");
        end

        266 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   266");
        end

        267 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   267");
        end

        268 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   268");
        end

        269 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   269");
        end

        270 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   270");
        end

        271 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   271");
        end

        272 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   272");
        end

        273 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   273");
        end

        274 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   274");
        end

        275 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   275");
        end

        276 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   276");
        end

        277 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   277");
        end

        278 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   278");
        end

        279 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   279");
        end

        280 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   280");
        end

        281 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   281");
        end

        282 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   282");
        end

        283 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   283");
        end

        284 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   284");
        end

        285 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   285");
        end

        286 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   286");
        end

        287 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   287");
        end

        288 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   288");
        end

        289 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   289");
        end

        290 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   290");
        end

        291 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   291");
        end

        292 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   292");
        end

        293 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   293");
        end

        294 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   294");
        end

        295 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   295");
        end

        296 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   296");
        end

        297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   297");
        end

        298 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   298");
        end

        299 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   299");
        end

        300 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   300");
        end

        301 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   301");
        end

        302 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   302");
        end

        303 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   303");
        end

        304 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   304");
        end

        305 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   305");
        end

        306 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   306");
        end

        307 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   307");
        end

        308 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   308");
        end

        309 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   309");
        end

        310 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   310");
        end

        311 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   311");
        end

        312 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   312");
        end

        313 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   313");
        end

        314 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   314");
        end

        315 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   315");
        end

        316 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   316");
        end

        317 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   317");
        end

        318 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   318");
        end

        319 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   319");
        end

        320 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   320");
        end

        321 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   321");
        end

        322 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   322");
        end

        323 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   323");
        end

        324 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   324");
        end

        325 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   325");
        end

        326 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   326");
        end

        327 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   327");
        end

        328 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   328");
        end

        329 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   329");
        end

        330 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   330");
        end

        331 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   331");
        end

        332 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   332");
        end

        333 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   333");
        end

        334 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   334");
        end

        335 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   335");
        end

        336 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   336");
        end

        337 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   337");
        end

        338 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   338");
        end

        339 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   339");
        end

        340 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   340");
        end

        341 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   341");
        end

        342 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   342");
        end

        343 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   343");
        end

        344 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   344");
        end

        345 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   345");
        end

        346 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   346");
        end

        347 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   347");
        end

        348 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   348");
        end

        349 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   349");
        end

        350 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   350");
        end

        351 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   351");
        end

        352 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   352");
        end

        353 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   353");
        end

        354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   354");
        end

        355 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   355");
        end

        356 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   356");
        end

        357 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   357");
        end

        358 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   358");
        end

        359 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   359");
        end

        360 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   360");
        end

        361 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   361");
        end

        362 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   362");
        end

        363 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   363");
        end

        364 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   364");
        end

        365 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   365");
        end

        366 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   366");
        end

        367 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   367");
        end

        368 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   368");
        end

        369 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   369");
        end

        370 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   370");
        end

        371 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   371");
        end

        372 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   372");
        end

        373 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   373");
        end

        374 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   374");
        end

        375 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   375");
        end

        376 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   376");
        end

        377 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   377");
        end

        378 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   378");
        end

        379 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   379");
        end

        380 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   380");
        end

        381 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   381");
        end

        382 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   382");
        end

        383 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   383");
        end

        384 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   384");
        end

        385 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   385");
        end

        386 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   386");
        end

        387 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   387");
        end

        388 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   388");
        end

        389 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   389");
        end

        390 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   390");
        end

        391 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   391");
        end

        392 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   392");
        end

        393 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   393");
        end

        394 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   394");
        end

        395 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   395");
        end

        396 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   396");
        end

        397 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   397");
        end

        398 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   398");
        end

        399 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   399");
        end

        400 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   400");
        end

        401 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   401");
        end

        402 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   402");
        end

        403 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   403");
        end

        404 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   404");
        end

        405 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   405");
        end

        406 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   406");
        end

        407 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   407");
        end

        408 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   408");
        end

        409 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   409");
        end

        410 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   410");
        end

        411 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   411");
        end

        412 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   412");
        end

        413 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   413");
        end

        414 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   414");
        end

        415 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   415");
        end

        416 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   416");
        end

        417 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   417");
        end

        418 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   418");
        end

        419 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   419");
        end

        420 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   420");
        end

        421 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   421");
        end

        422 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   422");
        end

        423 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   423");
        end

        424 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   424");
        end

        425 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   425");
        end

        426 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   426");
        end

        427 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   427");
        end

        428 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   428");
        end

        429 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   429");
        end

        430 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   430");
        end

        431 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   431");
        end

        432 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   432");
        end

        433 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   433");
        end

        434 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   434");
        end

        435 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   435");
        end

        436 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   436");
        end

        437 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   437");
        end

        438 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   438");
        end

        439 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   439");
        end

        440 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   440");
        end

        441 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   441");
        end

        442 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   442");
        end

        443 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   443");
        end

        444 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   444");
        end

        445 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   445");
        end

        446 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   446");
        end

        447 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   447");
        end

        448 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   448");
        end

        449 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   449");
        end

        450 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   450");
        end

        451 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   451");
        end

        452 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   452");
        end

        453 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   453");
        end

        454 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   454");
        end

        455 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   455");
        end

        456 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   456");
        end

        457 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   457");
        end

        458 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   458");
        end

        459 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   459");
        end

        460 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   460");
        end

        461 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   461");
        end

        462 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   462");
        end

        463 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   463");
        end

        464 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   464");
        end

        465 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   465");
        end

        466 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   466");
        end

        467 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   467");
        end

        468 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   468");
        end

        469 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   469");
        end

        470 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   470");
        end

        471 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   471");
        end

        472 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   472");
        end

        473 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   473");
        end

        474 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   474");
        end

        475 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   475");
        end

        476 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   476");
        end

        477 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   477");
        end

        478 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   478");
        end

        479 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   479");
        end

        480 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   480");
        end

        481 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   481");
        end

        482 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   482");
        end

        483 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   483");
        end

        484 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   484");
        end

        485 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   485");
        end

        486 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   486");
        end

        487 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   487");
        end

        488 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   488");
        end

        489 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   489");
        end

        490 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   490");
        end

        491 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   491");
        end

        492 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   492");
        end

        493 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   493");
        end

        494 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   494");
        end

        495 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   495");
        end

        496 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   496");
        end

        497 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   497");
        end

        498 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   498");
        end

        499 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   499");
        end

        500 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   500");
        end

        501 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   501");
        end

        502 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   502");
        end

        503 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   503");
        end

        504 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   504");
        end

        505 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   505");
        end

        506 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   506");
        end

        507 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   507");
        end

        508 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   508");
        end

        509 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   509");
        end

        510 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   510");
        end

        511 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   511");
        end

        512 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   512");
        end

        513 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   513");
        end

        514 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   514");
        end

        515 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   515");
        end

        516 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   516");
        end

        517 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   517");
        end

        518 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   518");
        end

        519 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   519");
        end

        520 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   520");
        end

        521 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   521");
        end

        522 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   522");
        end

        523 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   523");
        end

        524 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   524");
        end

        525 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   525");
        end

        526 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   526");
        end

        527 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   527");
        end

        528 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   528");
        end

        529 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   529");
        end

        530 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   530");
        end

        531 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   531");
        end

        532 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   532");
        end

        533 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   533");
        end

        534 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   534");
        end

        535 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   535");
        end

        536 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   536");
        end

        537 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   537");
        end

        538 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   538");
        end

        539 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   539");
        end

        540 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   540");
        end

        541 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   541");
        end

        542 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   542");
        end

        543 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   543");
        end

        544 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   544");
        end

        545 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   545");
        end

        546 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   546");
        end

        547 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   547");
        end

        548 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   548");
        end

        549 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   549");
        end

        550 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   550");
        end

        551 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   551");
        end

        552 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   552");
        end

        553 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   553");
        end

        554 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   554");
        end

        555 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   555");
        end

        556 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   556");
        end

        557 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   557");
        end

        558 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   558");
        end

        559 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   559");
        end

        560 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   560");
        end

        561 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   561");
        end

        562 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed   562");
        end

        563 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   563");
        end

        564 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   564");
        end

        565 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 566;
        end

        566 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 567;
              heapClock = 1;
        end

        567 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[81] = heapOut;
              ip = 568;
        end

        568 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 569;
        end

        569 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[619] = localMem[31];
              ip = 570;
        end

        570 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[619];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 571;
              heapClock = 1;
        end

        571 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 572;
        end

        572 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[620] = 0;
              ip = 573;
        end

        573 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[620];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 574;
              heapClock = 1;
        end

        574 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 575;
        end

        575 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 576;
              heapClock = 1;
        end

        576 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[82] = heapOut;
              ip = 577;
        end

        577 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 578;
        end

        578 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[621] = localMem[82];
              ip = 579;
        end

        579 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[621];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 580;
              heapClock = 1;
        end

        580 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 581;
        end

        581 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 582;
              heapClock = 1;
        end

        582 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[83] = heapOut;
              ip = 583;
        end

        583 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 584;
        end

        584 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[622] = localMem[83];
              ip = 585;
        end

        585 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[622];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 586;
              heapClock = 1;
        end

        586 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 587;
        end

        587 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[623] = 0;
              ip = 588;
        end

        588 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[623];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 589;
              heapClock = 1;
        end

        589 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 590;
        end

        590 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[624] = localMem[29];
              ip = 591;
        end

        591 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[624];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 592;
              heapClock = 1;
        end

        592 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 593;
        end

        593 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 594;
              heapClock = 1;
        end

        594 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 595;
        end

        595 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[625] = heapOut;                                                     // Data retrieved from heap memory
              ip = 596;
              heapClock = 1;
        end

        596 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 597;
        end

        597 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[626] = localMem[625] + 1;
              ip = 598;
        end

        598 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[29];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[626];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 599;
              heapClock = 1;
        end

        599 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 600;
        end

        600 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 601;
              heapClock = 1;
        end

        601 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 602;
        end

        602 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[627] = heapOut;                                                     // Data retrieved from heap memory
              ip = 603;
              heapClock = 1;
        end

        603 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 604;
        end

        604 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[628] = localMem[627];
              ip = 605;
        end

        605 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[628];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 606;
              heapClock = 1;
        end

        606 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 607;
        end

        607 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 608;
              heapClock = 1;
        end

        608 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[84] = heapOut;
              ip = 609;
        end

        609 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 610;
        end

        610 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[629] = localMem[31];
              ip = 611;
        end

        611 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[629];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 612;
              heapClock = 1;
        end

        612 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 613;
        end

        613 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[630] = 0;
              ip = 614;
        end

        614 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[630];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 615;
              heapClock = 1;
        end

        615 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 616;
        end

        616 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 617;
              heapClock = 1;
        end

        617 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[85] = heapOut;
              ip = 618;
        end

        618 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 619;
        end

        619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[631] = localMem[85];
              ip = 620;
        end

        620 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[631];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 621;
              heapClock = 1;
        end

        621 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 622;
        end

        622 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 623;
              heapClock = 1;
        end

        623 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[86] = heapOut;
              ip = 624;
        end

        624 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 625;
        end

        625 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[632] = localMem[86];
              ip = 626;
        end

        626 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[632];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 627;
              heapClock = 1;
        end

        627 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 628;
        end

        628 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[633] = 0;
              ip = 629;
        end

        629 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[633];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 630;
              heapClock = 1;
        end

        630 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 631;
        end

        631 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[634] = localMem[29];
              ip = 632;
        end

        632 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[634];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 633;
              heapClock = 1;
        end

        633 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 634;
        end

        634 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 635;
              heapClock = 1;
        end

        635 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 636;
        end

        636 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[635] = heapOut;                                                     // Data retrieved from heap memory
              ip = 637;
              heapClock = 1;
        end

        637 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 638;
        end

        638 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[636] = localMem[635] + 1;
              ip = 639;
        end

        639 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[29];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[636];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 640;
              heapClock = 1;
        end

        640 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 641;
        end

        641 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[29];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 642;
              heapClock = 1;
        end

        642 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 643;
        end

        643 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[637] = heapOut;                                                     // Data retrieved from heap memory
              ip = 644;
              heapClock = 1;
        end

        644 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 645;
        end

        645 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[638] = localMem[637];
              ip = 646;
        end

        646 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[638];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 647;
              heapClock = 1;
        end

        647 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 648;
        end

        648 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 649;
              heapClock = 1;
        end

        649 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 650;
        end

        650 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[639] = heapOut;                                                     // Data retrieved from heap memory
              ip = 651;
              heapClock = 1;
        end

        651 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 652;
        end

        652 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[87] = !localMem[639];
              ip = 653;
        end

        653 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[87] != 0 ? 795 : 654;
        end

        654 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 655;
              heapClock = 1;
        end

        655 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[88] = heapOut;
              ip = 656;
        end

        656 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 657;
        end

        657 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[640] = localMem[88];
              ip = 658;
        end

        658 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[640];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 659;
              heapClock = 1;
        end

        659 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 660;
        end

        660 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 661;
              heapClock = 1;
        end

        661 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[89] = heapOut;
              ip = 662;
        end

        662 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 663;
        end

        663 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[641] = localMem[89];
              ip = 664;
        end

        664 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[641];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 665;
              heapClock = 1;
        end

        665 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 666;
        end

        666 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 667;
              heapClock = 1;
        end

        667 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 668;
        end

        668 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[642] = heapOut;                                                     // Data retrieved from heap memory
              ip = 669;
              heapClock = 1;
        end

        669 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 670;
        end

        670 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[90] = localMem[642];
              ip = 671;
        end

        671 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 672;
              heapClock = 1;
        end

        672 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 673;
        end

        673 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[643] = heapOut;                                                     // Data retrieved from heap memory
              ip = 674;
              heapClock = 1;
        end

        674 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 675;
        end

        675 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[91] = localMem[643];
              ip = 676;
        end

        676 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[90];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 677;
              heapClock = 1;
        end

        677 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[91];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 678;
              heapClock = 1;
        end

        678 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 679;
              heapClock = 1;
        end

        679 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 680;
        end

        680 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[644] = heapOut;                                                     // Data retrieved from heap memory
              ip = 681;
              heapClock = 1;
        end

        681 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 682;
        end

        682 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[92] = localMem[644];
              ip = 683;
        end

        683 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 684;
              heapClock = 1;
        end

        684 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 685;
        end

        685 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[645] = heapOut;                                                     // Data retrieved from heap memory
              ip = 686;
              heapClock = 1;
        end

        686 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 687;
        end

        687 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[93] = localMem[645];
              ip = 688;
        end

        688 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[92];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 689;
              heapClock = 1;
        end

        689 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[93];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 690;
              heapClock = 1;
        end

        690 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 691;
              heapClock = 1;
        end

        691 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 692;
        end

        692 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[646] = heapOut;                                                     // Data retrieved from heap memory
              ip = 693;
              heapClock = 1;
        end

        693 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 694;
        end

        694 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[94] = localMem[646];
              ip = 695;
        end

        695 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 696;
              heapClock = 1;
        end

        696 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 697;
        end

        697 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[647] = heapOut;                                                     // Data retrieved from heap memory
              ip = 698;
              heapClock = 1;
        end

        698 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 699;
        end

        699 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[95] = localMem[647];
              ip = 700;
        end

        700 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[96] = localMem[31] + 1;
              ip = 701;
        end

        701 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[94];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 702;
              heapClock = 1;
        end

        702 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[95];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[96];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 703;
              heapClock = 1;
        end

        703 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 704;
              heapClock = 1;
        end

        704 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 705;
        end

        705 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[648] = heapOut;                                                     // Data retrieved from heap memory
              ip = 706;
              heapClock = 1;
        end

        706 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 707;
        end

        707 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[97] = localMem[648];
              ip = 708;
        end

        708 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 709;
              heapClock = 1;
        end

        709 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 710;
        end

        710 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[649] = heapOut;                                                     // Data retrieved from heap memory
              ip = 711;
              heapClock = 1;
        end

        711 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 712;
        end

        712 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[98] = localMem[649];
              ip = 713;
        end

        713 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[97];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 714;
              heapClock = 1;
        end

        714 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[98];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 715;
              heapClock = 1;
        end

        715 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 716;
              heapClock = 1;
        end

        716 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 717;
        end

        717 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[650] = heapOut;                                                     // Data retrieved from heap memory
              ip = 718;
              heapClock = 1;
        end

        718 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 719;
        end

        719 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[99] = localMem[650];
              ip = 720;
        end

        720 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 721;
              heapClock = 1;
        end

        721 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 722;
        end

        722 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[651] = heapOut;                                                     // Data retrieved from heap memory
              ip = 723;
              heapClock = 1;
        end

        723 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 724;
        end

        724 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[100] = localMem[651];
              ip = 725;
        end

        725 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[99];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 726;
              heapClock = 1;
        end

        726 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[100];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 727;
              heapClock = 1;
        end

        727 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 728;
              heapClock = 1;
        end

        728 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 729;
        end

        729 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[652] = heapOut;                                                     // Data retrieved from heap memory
              ip = 730;
              heapClock = 1;
        end

        730 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 731;
        end

        731 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[101] = localMem[652];
              ip = 732;
        end

        732 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 733;
              heapClock = 1;
        end

        733 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 734;
        end

        734 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[653] = heapOut;                                                     // Data retrieved from heap memory
              ip = 735;
              heapClock = 1;
        end

        735 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 736;
        end

        736 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[102] = localMem[653];
              ip = 737;
        end

        737 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[103] = localMem[31] + 1;
              ip = 738;
        end

        738 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[101];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 739;
              heapClock = 1;
        end

        739 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[102];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[103];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 740;
              heapClock = 1;
        end

        740 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 741;
              heapClock = 1;
        end

        741 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 742;
        end

        742 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[654] = heapOut;                                                     // Data retrieved from heap memory
              ip = 743;
              heapClock = 1;
        end

        743 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 744;
        end

        744 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[104] = localMem[654];
              ip = 745;
        end

        745 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[105] = localMem[104] + 1;
              ip = 746;
        end

        746 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 747;
              heapClock = 1;
        end

        747 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 748;
        end

        748 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[655] = heapOut;                                                     // Data retrieved from heap memory
              ip = 749;
              heapClock = 1;
        end

        749 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 750;
        end

        750 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[106] = localMem[655];
              ip = 751;
        end

        751 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 752;
        end

        752 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[107] = 0;
              ip = 753;
        end

        753 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 754;
        end

        754 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[107] >= localMem[105] ? 766 : 755;
        end

        755 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[106];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[107];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 756;
              heapClock = 1;
        end

        756 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 757;
        end

        757 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[656] = heapOut;                                                     // Data retrieved from heap memory
              ip = 758;
              heapClock = 1;
        end

        758 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 759;
        end

        759 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[108] = localMem[656];
              ip = 760;
        end

        760 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[657] = localMem[81];
              ip = 761;
        end

        761 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[108];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[657];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 762;
              heapClock = 1;
        end

        762 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 763;
        end

        763 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 764;
        end

        764 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[107] = localMem[107] + 1;
              ip = 765;
        end

        765 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 753;
        end

        766 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 767;
        end

        767 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 768;
              heapClock = 1;
        end

        768 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 769;
        end

        769 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[658] = heapOut;                                                     // Data retrieved from heap memory
              ip = 770;
              heapClock = 1;
        end

        770 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 771;
        end

        771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[109] = localMem[658];
              ip = 772;
        end

        772 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[110] = localMem[109] + 1;
              ip = 773;
        end

        773 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 774;
              heapClock = 1;
        end

        774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 775;
        end

        775 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[659] = heapOut;                                                     // Data retrieved from heap memory
              ip = 776;
              heapClock = 1;
        end

        776 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 777;
        end

        777 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[111] = localMem[659];
              ip = 778;
        end

        778 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 779;
        end

        779 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[112] = 0;
              ip = 780;
        end

        780 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 781;
        end

        781 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[112] >= localMem[110] ? 793 : 782;
        end

        782 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[111];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[112];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 783;
              heapClock = 1;
        end

        783 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 784;
        end

        784 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[660] = heapOut;                                                     // Data retrieved from heap memory
              ip = 785;
              heapClock = 1;
        end

        785 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 786;
        end

        786 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[113] = localMem[660];
              ip = 787;
        end

        787 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[661] = localMem[84];
              ip = 788;
        end

        788 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[113];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[661];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 789;
              heapClock = 1;
        end

        789 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 790;
        end

        790 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 791;
        end

        791 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[112] = localMem[112] + 1;
              ip = 792;
        end

        792 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 780;
        end

        793 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 794;
        end

        794 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 850;
        end

        795 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 796;
        end

        796 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 797;
              heapClock = 1;
        end

        797 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[114] = heapOut;
              ip = 798;
        end

        798 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 799;
        end

        799 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[662] = localMem[114];
              ip = 800;
        end

        800 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[26];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[662];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 801;
              heapClock = 1;
        end

        801 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 802;
        end

        802 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 803;
              heapClock = 1;
        end

        803 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 804;
        end

        804 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[663] = heapOut;                                                     // Data retrieved from heap memory
              ip = 805;
              heapClock = 1;
        end

        805 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 806;
        end

        806 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[115] = localMem[663];
              ip = 807;
        end

        807 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 808;
              heapClock = 1;
        end

        808 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 809;
        end

        809 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[664] = heapOut;                                                     // Data retrieved from heap memory
              ip = 810;
              heapClock = 1;
        end

        810 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 811;
        end

        811 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[116] = localMem[664];
              ip = 812;
        end

        812 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[115];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 813;
              heapClock = 1;
        end

        813 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[116];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 814;
              heapClock = 1;
        end

        814 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 815;
              heapClock = 1;
        end

        815 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 816;
        end

        816 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[665] = heapOut;                                                     // Data retrieved from heap memory
              ip = 817;
              heapClock = 1;
        end

        817 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 818;
        end

        818 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[117] = localMem[665];
              ip = 819;
        end

        819 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[81];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 820;
              heapClock = 1;
        end

        820 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 821;
        end

        821 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[666] = heapOut;                                                     // Data retrieved from heap memory
              ip = 822;
              heapClock = 1;
        end

        822 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 823;
        end

        823 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[118] = localMem[666];
              ip = 824;
        end

        824 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[117];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 825;
              heapClock = 1;
        end

        825 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[118];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 826;
              heapClock = 1;
        end

        826 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 827;
              heapClock = 1;
        end

        827 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 828;
        end

        828 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[667] = heapOut;                                                     // Data retrieved from heap memory
              ip = 829;
              heapClock = 1;
        end

        829 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 830;
        end

        830 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[119] = localMem[667];
              ip = 831;
        end

        831 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 832;
              heapClock = 1;
        end

        832 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 833;
        end

        833 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[668] = heapOut;                                                     // Data retrieved from heap memory
              ip = 834;
              heapClock = 1;
        end

        834 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 835;
        end

        835 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[120] = localMem[668];
              ip = 836;
        end

        836 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[119];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 837;
              heapClock = 1;
        end

        837 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[120];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 838;
              heapClock = 1;
        end

        838 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 839;
              heapClock = 1;
        end

        839 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 840;
        end

        840 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[669] = heapOut;                                                     // Data retrieved from heap memory
              ip = 841;
              heapClock = 1;
        end

        841 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 842;
        end

        842 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[121] = localMem[669];
              ip = 843;
        end

        843 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[84];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 844;
              heapClock = 1;
        end

        844 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 845;
        end

        845 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[670] = heapOut;                                                     // Data retrieved from heap memory
              ip = 846;
              heapClock = 1;
        end

        846 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 847;
        end

        847 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[122] = localMem[670];
              ip = 848;
        end

        848 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[121];                                                 // Array to write to
              heapIndex  = localMem[32];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 849;
              heapClock = 1;
        end

        849 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[122];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[31];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 850;
              heapClock = 1;
        end

        850 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 851;
        end

        851 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[671] = localMem[26];
              ip = 852;
        end

        852 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[81];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[671];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 853;
              heapClock = 1;
        end

        853 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 854;
        end

        854 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[672] = localMem[26];
              ip = 855;
        end

        855 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[84];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[672];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 856;
              heapClock = 1;
        end

        856 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 857;
        end

        857 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 858;
              heapClock = 1;
        end

        858 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 859;
        end

        859 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[673] = heapOut;                                                     // Data retrieved from heap memory
              ip = 860;
              heapClock = 1;
        end

        860 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 861;
        end

        861 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[123] = localMem[673];
              ip = 862;
        end

        862 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[123];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 863;
              heapClock = 1;
        end

        863 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 864;
        end

        864 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[674] = heapOut;                                                     // Data retrieved from heap memory
              ip = 865;
              heapClock = 1;
        end

        865 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 866;
        end

        866 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[124] = localMem[674];
              ip = 867;
        end

        867 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 868;
              heapClock = 1;
        end

        868 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 869;
        end

        869 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[675] = heapOut;                                                     // Data retrieved from heap memory
              ip = 870;
              heapClock = 1;
        end

        870 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 871;
        end

        871 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[125] = localMem[675];
              ip = 872;
        end

        872 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[125];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 873;
              heapClock = 1;
        end

        873 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 874;
        end

        874 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[676] = heapOut;                                                     // Data retrieved from heap memory
              ip = 875;
              heapClock = 1;
        end

        875 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 876;
        end

        876 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[126] = localMem[676];
              ip = 877;
        end

        877 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 878;
              heapClock = 1;
        end

        878 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 879;
        end

        879 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[677] = heapOut;                                                     // Data retrieved from heap memory
              ip = 880;
              heapClock = 1;
        end

        880 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 881;
        end

        881 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[127] = localMem[677];
              ip = 882;
        end

        882 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[678] = localMem[124];
              ip = 883;
        end

        883 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[127];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[678];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 884;
              heapClock = 1;
        end

        884 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 885;
        end

        885 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 886;
              heapClock = 1;
        end

        886 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 887;
        end

        887 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[679] = heapOut;                                                     // Data retrieved from heap memory
              ip = 888;
              heapClock = 1;
        end

        888 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 889;
        end

        889 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[128] = localMem[679];
              ip = 890;
        end

        890 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[680] = localMem[126];
              ip = 891;
        end

        891 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[128];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[680];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 892;
              heapClock = 1;
        end

        892 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 893;
        end

        893 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 894;
              heapClock = 1;
        end

        894 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 895;
        end

        895 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[681] = heapOut;                                                     // Data retrieved from heap memory
              ip = 896;
              heapClock = 1;
        end

        896 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 897;
        end

        897 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[129] = localMem[681];
              ip = 898;
        end

        898 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[682] = localMem[81];
              ip = 899;
        end

        899 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[129];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[682];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 900;
              heapClock = 1;
        end

        900 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 901;
        end

        901 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 902;
              heapClock = 1;
        end

        902 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 903;
        end

        903 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[683] = heapOut;                                                     // Data retrieved from heap memory
              ip = 904;
              heapClock = 1;
        end

        904 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 905;
        end

        905 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[130] = localMem[683];
              ip = 906;
        end

        906 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[684] = localMem[84];
              ip = 907;
        end

        907 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[130];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[684];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 908;
              heapClock = 1;
        end

        908 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 909;
        end

        909 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[685] = 1;
              ip = 910;
        end

        910 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[26];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[685];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 911;
              heapClock = 1;
        end

        911 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 912;
        end

        912 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 913;
              heapClock = 1;
        end

        913 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 914;
        end

        914 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[686] = heapOut;                                                     // Data retrieved from heap memory
              ip = 915;
              heapClock = 1;
        end

        915 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 916;
        end

        916 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[131] = localMem[686];
              ip = 917;
        end

        917 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[131];
              ip = 918;
              heapClock = 1;
        end

        918 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 919;
              heapClock = 1;
        end

        919 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 920;
        end

        920 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[687] = heapOut;                                                     // Data retrieved from heap memory
              ip = 921;
              heapClock = 1;
        end

        921 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 922;
        end

        922 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[132] = localMem[687];
              ip = 923;
        end

        923 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[132];
              ip = 924;
              heapClock = 1;
        end

        924 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 925;
              heapClock = 1;
        end

        925 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 926;
        end

        926 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[688] = heapOut;                                                     // Data retrieved from heap memory
              ip = 927;
              heapClock = 1;
        end

        927 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 928;
        end

        928 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[133] = localMem[688];
              ip = 929;
        end

        929 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 2;
              heapArray  = localMem[133];
              ip = 930;
              heapClock = 1;
        end

        930 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 932;
        end

        931 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   931");
        end

        932 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 933;
        end

        933 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[27] = 1;
              ip = 934;
        end

        934 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 937;
        end

        935 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 936;
        end

        936 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[27] = 0;
              ip = 937;
        end

        937 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 938;
        end

        938 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 939;
        end

        939 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 940;
        end

        940 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[134] = 0;
              ip = 941;
        end

        941 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 942;
        end

        942 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[134] >= 99 ? 2456 : 943;
        end

        943 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 944;
              heapClock = 1;
        end

        944 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 945;
        end

        945 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[689] = heapOut;                                                     // Data retrieved from heap memory
              ip = 946;
              heapClock = 1;
        end

        946 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 947;
        end

        947 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[135] = localMem[689];
              ip = 948;
        end

        948 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[136] = localMem[135] - 1;
              ip = 949;
        end

        949 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 950;
              heapClock = 1;
        end

        950 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 951;
        end

        951 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[690] = heapOut;                                                     // Data retrieved from heap memory
              ip = 952;
              heapClock = 1;
        end

        952 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 953;
        end

        953 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[137] = localMem[690];
              ip = 954;
        end

        954 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[137];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[136];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 955;
              heapClock = 1;
        end

        955 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 956;
        end

        956 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[691] = heapOut;                                                     // Data retrieved from heap memory
              ip = 957;
              heapClock = 1;
        end

        957 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 958;
        end

        958 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[138] = localMem[691];
              ip = 959;
        end

        959 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[1] <= localMem[138] ? 1695 : 960;
        end

        960 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 961;
              heapClock = 1;
        end

        961 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 962;
        end

        962 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[692] = heapOut;                                                     // Data retrieved from heap memory
              ip = 963;
              heapClock = 1;
        end

        963 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 964;
        end

        964 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[139] = !localMem[692];
              ip = 965;
        end

        965 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[139] == 0 ? 976 : 966;
        end

        966 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[693] = localMem[26];
              ip = 967;
        end

        967 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[693];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 968;
              heapClock = 1;
        end

        968 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 969;
        end

        969 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[694] = 2;
              ip = 970;
        end

        970 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[694];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 971;
              heapClock = 1;
        end

        971 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 972;
        end

        972 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[695] = localMem[135] - 1;
              ip = 973;
        end

        973 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[695];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 974;
              heapClock = 1;
        end

        974 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 975;
        end

        975 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2460;
        end

        976 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 977;
        end

        977 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[26];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 978;
              heapClock = 1;
        end

        978 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 979;
        end

        979 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[696] = heapOut;                                                     // Data retrieved from heap memory
              ip = 980;
              heapClock = 1;
        end

        980 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 981;
        end

        981 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[140] = localMem[696];
              ip = 982;
        end

        982 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[135];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 983;
              heapClock = 1;
        end

        983 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 984;
        end

        984 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[697] = heapOut;                                                     // Data retrieved from heap memory
              ip = 985;
              heapClock = 1;
        end

        985 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 986;
        end

        986 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[141] = localMem[697];
              ip = 987;
        end

        987 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 988;
        end

        988 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 989;
              heapClock = 1;
        end

        989 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 990;
        end

        990 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[698] = heapOut;                                                     // Data retrieved from heap memory
              ip = 991;
              heapClock = 1;
        end

        991 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 992;
        end

        992 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[143] = localMem[698];
              ip = 993;
        end

        993 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 994;
              heapClock = 1;
        end

        994 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 995;
        end

        995 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[699] = heapOut;                                                     // Data retrieved from heap memory
              ip = 996;
              heapClock = 1;
        end

        996 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 997;
        end

        997 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[144] = localMem[699];
              ip = 998;
        end

        998 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 999;
              heapClock = 1;
        end

        999 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1000;
        end

       1000 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[700] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1001;
              heapClock = 1;
        end

       1001 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1002;
        end

       1002 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[145] = localMem[700];
              ip = 1003;
        end

       1003 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[143] <  localMem[145] ? 1688 : 1004;
        end

       1004 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[146] = localMem[145];
              ip = 1005;
        end

       1005 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[146] = localMem[146] >> 1;
              ip = 1006;
              ip = 1006;
        end

       1006 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[147] = localMem[146] + 1;
              ip = 1007;
        end

       1007 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1008;
              heapClock = 1;
        end

       1008 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1009;
        end

       1009 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[701] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1010;
              heapClock = 1;
        end

       1010 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1011;
        end

       1011 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[148] = localMem[701];
              ip = 1012;
        end

       1012 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[148] == 0 ? 1318 : 1013;
        end

       1013 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1014;
              heapClock = 1;
        end

       1014 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[149] = heapOut;
              ip = 1015;
        end

       1015 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1016;
        end

       1016 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[702] = localMem[146];
              ip = 1017;
        end

       1017 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[702];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1018;
              heapClock = 1;
        end

       1018 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1019;
        end

       1019 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[703] = 0;
              ip = 1020;
        end

       1020 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[703];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1021;
              heapClock = 1;
        end

       1021 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1022;
        end

       1022 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1023;
              heapClock = 1;
        end

       1023 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[150] = heapOut;
              ip = 1024;
        end

       1024 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1025;
        end

       1025 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[704] = localMem[150];
              ip = 1026;
        end

       1026 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[704];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1027;
              heapClock = 1;
        end

       1027 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1028;
        end

       1028 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1029;
              heapClock = 1;
        end

       1029 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[151] = heapOut;
              ip = 1030;
        end

       1030 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1031;
        end

       1031 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[705] = localMem[151];
              ip = 1032;
        end

       1032 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[705];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1033;
              heapClock = 1;
        end

       1033 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1034;
        end

       1034 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[706] = 0;
              ip = 1035;
        end

       1035 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[706];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1036;
              heapClock = 1;
        end

       1036 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1037;
        end

       1037 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[707] = localMem[144];
              ip = 1038;
        end

       1038 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[707];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1039;
              heapClock = 1;
        end

       1039 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1040;
        end

       1040 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1041;
              heapClock = 1;
        end

       1041 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1042;
        end

       1042 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[708] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1043;
              heapClock = 1;
        end

       1043 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1044;
        end

       1044 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[709] = localMem[708] + 1;
              ip = 1045;
        end

       1045 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[144];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[709];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1046;
              heapClock = 1;
        end

       1046 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1047;
        end

       1047 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1048;
              heapClock = 1;
        end

       1048 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1049;
        end

       1049 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[710] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1050;
              heapClock = 1;
        end

       1050 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1051;
        end

       1051 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[711] = localMem[710];
              ip = 1052;
        end

       1052 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[711];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1053;
              heapClock = 1;
        end

       1053 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1054;
        end

       1054 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1055;
              heapClock = 1;
        end

       1055 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1056;
        end

       1056 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[712] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1057;
              heapClock = 1;
        end

       1057 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1058;
        end

       1058 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[152] = !localMem[712];
              ip = 1059;
        end

       1059 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[152] != 0 ? 1137 : 1060;
        end

       1060 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1061;
              heapClock = 1;
        end

       1061 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[153] = heapOut;
              ip = 1062;
        end

       1062 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1063;
        end

       1063 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[713] = localMem[153];
              ip = 1064;
        end

       1064 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[713];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1065;
              heapClock = 1;
        end

       1065 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1066;
        end

       1066 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1067;
              heapClock = 1;
        end

       1067 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1068;
        end

       1068 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[714] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1069;
              heapClock = 1;
        end

       1069 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1070;
        end

       1070 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[154] = localMem[714];
              ip = 1071;
        end

       1071 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1072;
              heapClock = 1;
        end

       1072 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1073;
        end

       1073 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[715] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1074;
              heapClock = 1;
        end

       1074 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1075;
        end

       1075 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[155] = localMem[715];
              ip = 1076;
        end

       1076 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[154];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1077;
              heapClock = 1;
        end

       1077 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[155];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[146];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1078;
              heapClock = 1;
        end

       1078 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1079;
              heapClock = 1;
        end

       1079 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1080;
        end

       1080 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[716] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1081;
              heapClock = 1;
        end

       1081 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1082;
        end

       1082 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[156] = localMem[716];
              ip = 1083;
        end

       1083 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1084;
              heapClock = 1;
        end

       1084 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1085;
        end

       1085 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[717] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1086;
              heapClock = 1;
        end

       1086 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1087;
        end

       1087 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[157] = localMem[717];
              ip = 1088;
        end

       1088 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[156];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1089;
              heapClock = 1;
        end

       1089 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[157];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[146];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1090;
              heapClock = 1;
        end

       1090 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1091;
              heapClock = 1;
        end

       1091 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1092;
        end

       1092 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[718] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1093;
              heapClock = 1;
        end

       1093 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1094;
        end

       1094 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[158] = localMem[718];
              ip = 1095;
        end

       1095 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1096;
              heapClock = 1;
        end

       1096 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1097;
        end

       1097 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[719] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1098;
              heapClock = 1;
        end

       1098 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1099;
        end

       1099 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[159] = localMem[719];
              ip = 1100;
        end

       1100 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[160] = localMem[146] + 1;
              ip = 1101;
        end

       1101 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[158];                                                 // Array to write to
              heapIndex  = localMem[147];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1102;
              heapClock = 1;
        end

       1102 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[159];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[160];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1103;
              heapClock = 1;
        end

       1103 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1104;
              heapClock = 1;
        end

       1104 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1105;
        end

       1105 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[720] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1106;
              heapClock = 1;
        end

       1106 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1107;
        end

       1107 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[161] = localMem[720];
              ip = 1108;
        end

       1108 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[162] = localMem[161] + 1;
              ip = 1109;
        end

       1109 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[149];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1110;
              heapClock = 1;
        end

       1110 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1111;
        end

       1111 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[721] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1112;
              heapClock = 1;
        end

       1112 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1113;
        end

       1113 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[163] = localMem[721];
              ip = 1114;
        end

       1114 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1115;
        end

       1115 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[164] = 0;
              ip = 1116;
        end

       1116 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1117;
        end

       1117 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[164] >= localMem[162] ? 1129 : 1118;
        end

       1118 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[163];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[164];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1119;
              heapClock = 1;
        end

       1119 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1120;
        end

       1120 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[722] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1121;
              heapClock = 1;
        end

       1121 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1122;
        end

       1122 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[165] = localMem[722];
              ip = 1123;
        end

       1123 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[723] = localMem[149];
              ip = 1124;
        end

       1124 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[165];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[723];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1125;
              heapClock = 1;
        end

       1125 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1126;
        end

       1126 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1127;
        end

       1127 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[164] = localMem[164] + 1;
              ip = 1128;
        end

       1128 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1116;
        end

       1129 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1130;
        end

       1130 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1131;
              heapClock = 1;
        end

       1131 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1132;
        end

       1132 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[724] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1133;
              heapClock = 1;
        end

       1133 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1134;
        end

       1134 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[166] = localMem[724];
              ip = 1135;
        end

       1135 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[147];
              heapArray  = localMem[166];
              ip = 1136;
              heapClock = 1;
        end

       1136 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1162;
        end

       1137 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1137");
        end

       1138 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1138");
        end

       1139 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1139");
        end

       1140 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1140");
        end

       1141 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1141");
        end

       1142 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1142");
        end

       1143 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1143");
        end

       1144 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1144");
        end

       1145 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1145");
        end

       1146 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1146");
        end

       1147 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1147");
        end

       1148 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1148");
        end

       1149 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1149");
        end

       1150 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1150");
        end

       1151 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1151");
        end

       1152 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1152");
        end

       1153 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1153");
        end

       1154 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1154");
        end

       1155 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1155");
        end

       1156 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1156");
        end

       1157 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1157");
        end

       1158 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1158");
        end

       1159 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1159");
        end

       1160 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1160");
        end

       1161 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1161");
        end

       1162 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1163;
        end

       1163 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[729] = localMem[146];
              ip = 1164;
        end

       1164 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[141];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[729];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1165;
              heapClock = 1;
        end

       1165 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1166;
        end

       1166 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[730] = localMem[148];
              ip = 1167;
        end

       1167 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[149];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[730];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1168;
              heapClock = 1;
        end

       1168 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1169;
        end

       1169 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1170;
              heapClock = 1;
        end

       1170 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1171;
        end

       1171 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[731] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1172;
              heapClock = 1;
        end

       1172 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1173;
        end

       1173 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[171] = localMem[731];
              ip = 1174;
        end

       1174 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1175;
              heapClock = 1;
        end

       1175 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1176;
        end

       1176 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[732] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1177;
              heapClock = 1;
        end

       1177 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1178;
        end

       1178 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[172] = localMem[732];
              ip = 1179;
        end

       1179 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[172];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[171];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1180;
              heapClock = 1;
        end

       1180 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1181;
        end

       1181 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[733] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1182;
              heapClock = 1;
        end

       1182 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1183;
        end

       1183 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[173] = localMem[733];
              ip = 1184;
        end

       1184 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[173] != localMem[141] ? 1247 : 1185;
        end

       1185 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1186;
              heapClock = 1;
        end

       1186 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1187;
        end

       1187 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[734] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1188;
              heapClock = 1;
        end

       1188 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1189;
        end

       1189 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[174] = localMem[734];
              ip = 1190;
        end

       1190 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[174];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[146];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1191;
              heapClock = 1;
        end

       1191 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1192;
        end

       1192 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[735] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1193;
              heapClock = 1;
        end

       1193 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1194;
        end

       1194 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[175] = localMem[735];
              ip = 1195;
        end

       1195 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1196;
              heapClock = 1;
        end

       1196 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1197;
        end

       1197 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[736] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1198;
              heapClock = 1;
        end

       1198 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1199;
        end

       1199 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[176] = localMem[736];
              ip = 1200;
        end

       1200 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[737] = localMem[175];
              ip = 1201;
        end

       1201 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[176];                                                // Array to write to
              heapIndex   = localMem[171];                                                // Index of element to write to
              heapIn      = localMem[737];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1202;
              heapClock = 1;
        end

       1202 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1203;
        end

       1203 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1204;
              heapClock = 1;
        end

       1204 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1205;
        end

       1205 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[738] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1206;
              heapClock = 1;
        end

       1206 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1207;
        end

       1207 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[177] = localMem[738];
              ip = 1208;
        end

       1208 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[177];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[146];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1209;
              heapClock = 1;
        end

       1209 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1210;
        end

       1210 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[739] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1211;
              heapClock = 1;
        end

       1211 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1212;
        end

       1212 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[178] = localMem[739];
              ip = 1213;
        end

       1213 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1214;
              heapClock = 1;
        end

       1214 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1215;
        end

       1215 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[740] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1216;
              heapClock = 1;
        end

       1216 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1217;
        end

       1217 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[179] = localMem[740];
              ip = 1218;
        end

       1218 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[741] = localMem[178];
              ip = 1219;
        end

       1219 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[179];                                                // Array to write to
              heapIndex   = localMem[171];                                                // Index of element to write to
              heapIn      = localMem[741];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1220;
              heapClock = 1;
        end

       1220 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1221;
        end

       1221 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1222;
              heapClock = 1;
        end

       1222 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1223;
        end

       1223 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[742] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1224;
              heapClock = 1;
        end

       1224 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1225;
        end

       1225 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[180] = localMem[742];
              ip = 1226;
        end

       1226 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[146];
              heapArray  = localMem[180];
              ip = 1227;
              heapClock = 1;
        end

       1227 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[141];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1228;
              heapClock = 1;
        end

       1228 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1229;
        end

       1229 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[743] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1230;
              heapClock = 1;
        end

       1230 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1231;
        end

       1231 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[181] = localMem[743];
              ip = 1232;
        end

       1232 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[146];
              heapArray  = localMem[181];
              ip = 1233;
              heapClock = 1;
        end

       1233 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[182] = localMem[171] + 1;
              ip = 1234;
        end

       1234 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[744] = localMem[182];
              ip = 1235;
        end

       1235 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[148];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[744];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1236;
              heapClock = 1;
        end

       1236 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1237;
        end

       1237 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[148];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1238;
              heapClock = 1;
        end

       1238 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1239;
        end

       1239 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[745] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1240;
              heapClock = 1;
        end

       1240 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1241;
        end

       1241 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[183] = localMem[745];
              ip = 1242;
        end

       1242 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[746] = localMem[149];
              ip = 1243;
        end

       1243 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[183];                                                // Array to write to
              heapIndex   = localMem[182];                                                // Index of element to write to
              heapIn      = localMem[746];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1244;
              heapClock = 1;
        end

       1244 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 1245;
        end

       1245 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1685;
        end

       1246 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1246");
        end

       1247 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1247");
        end

       1248 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  1248");
        end

       1249 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1249");
        end

       1250 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1250");
        end

       1251 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1251");
        end

       1252 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1252");
        end

       1253 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1253");
        end

       1254 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1254");
        end

       1255 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1255");
        end

       1256 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1256");
        end

       1257 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1257");
        end

       1258 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1258");
        end

       1259 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1259");
        end

       1260 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1260");
        end

       1261 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1261");
        end

       1262 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1262");
        end

       1263 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1263");
        end

       1264 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1264");
        end

       1265 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1265");
        end

       1266 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1266");
        end

       1267 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1267");
        end

       1268 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1268");
        end

       1269 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1269");
        end

       1270 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1270");
        end

       1271 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1271");
        end

       1272 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1272");
        end

       1273 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1273");
        end

       1274 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1274");
        end

       1275 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1275");
        end

       1276 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1276");
        end

       1277 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1277");
        end

       1278 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1278");
        end

       1279 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1279");
        end

       1280 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1280");
        end

       1281 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1281");
        end

       1282 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1282");
        end

       1283 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1283");
        end

       1284 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1284");
        end

       1285 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1285");
        end

       1286 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1286");
        end

       1287 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1287");
        end

       1288 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1288");
        end

       1289 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1289");
        end

       1290 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1290");
        end

       1291 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1291");
        end

       1292 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1292");
        end

       1293 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1293");
        end

       1294 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1294");
        end

       1295 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1295");
        end

       1296 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1296");
        end

       1297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1297");
        end

       1298 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1298");
        end

       1299 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1299");
        end

       1300 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1300");
        end

       1301 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1301");
        end

       1302 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1302");
        end

       1303 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1303");
        end

       1304 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1304");
        end

       1305 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1305");
        end

       1306 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1306");
        end

       1307 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1307");
        end

       1308 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1308");
        end

       1309 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1309");
        end

       1310 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1310");
        end

       1311 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1311");
        end

       1312 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1312");
        end

       1313 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1313");
        end

       1314 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1314");
        end

       1315 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1315");
        end

       1316 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1316");
        end

       1317 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1317");
        end

       1318 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1318");
        end

       1319 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1319");
        end

       1320 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1320");
        end

       1321 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1321");
        end

       1322 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1322");
        end

       1323 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1323");
        end

       1324 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1324");
        end

       1325 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1325");
        end

       1326 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1326");
        end

       1327 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1327");
        end

       1328 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1328");
        end

       1329 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1329");
        end

       1330 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1330");
        end

       1331 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1331");
        end

       1332 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1332");
        end

       1333 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1333");
        end

       1334 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1334");
        end

       1335 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1335");
        end

       1336 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1336");
        end

       1337 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1337");
        end

       1338 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1338");
        end

       1339 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1339");
        end

       1340 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1340");
        end

       1341 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1341");
        end

       1342 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1342");
        end

       1343 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1343");
        end

       1344 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1344");
        end

       1345 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1345");
        end

       1346 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1346");
        end

       1347 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1347");
        end

       1348 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1348");
        end

       1349 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1349");
        end

       1350 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1350");
        end

       1351 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1351");
        end

       1352 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1352");
        end

       1353 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1353");
        end

       1354 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1354");
        end

       1355 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1355");
        end

       1356 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1356");
        end

       1357 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1357");
        end

       1358 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1358");
        end

       1359 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1359");
        end

       1360 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1360");
        end

       1361 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1361");
        end

       1362 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1362");
        end

       1363 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1363");
        end

       1364 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1364");
        end

       1365 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1365");
        end

       1366 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1366");
        end

       1367 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1367");
        end

       1368 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1368");
        end

       1369 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1369");
        end

       1370 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1370");
        end

       1371 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1371");
        end

       1372 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1372");
        end

       1373 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1373");
        end

       1374 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1374");
        end

       1375 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1375");
        end

       1376 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1376");
        end

       1377 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1377");
        end

       1378 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1378");
        end

       1379 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1379");
        end

       1380 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1380");
        end

       1381 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1381");
        end

       1382 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1382");
        end

       1383 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1383");
        end

       1384 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1384");
        end

       1385 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1385");
        end

       1386 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1386");
        end

       1387 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1387");
        end

       1388 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1388");
        end

       1389 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1389");
        end

       1390 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1390");
        end

       1391 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1391");
        end

       1392 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1392");
        end

       1393 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1393");
        end

       1394 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1394");
        end

       1395 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1395");
        end

       1396 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1396");
        end

       1397 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1397");
        end

       1398 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1398");
        end

       1399 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1399");
        end

       1400 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1400");
        end

       1401 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1401");
        end

       1402 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1402");
        end

       1403 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1403");
        end

       1404 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1404");
        end

       1405 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1405");
        end

       1406 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1406");
        end

       1407 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1407");
        end

       1408 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1408");
        end

       1409 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1409");
        end

       1410 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1410");
        end

       1411 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1411");
        end

       1412 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1412");
        end

       1413 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1413");
        end

       1414 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1414");
        end

       1415 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1415");
        end

       1416 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1416");
        end

       1417 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1417");
        end

       1418 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1418");
        end

       1419 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1419");
        end

       1420 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1420");
        end

       1421 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1421");
        end

       1422 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1422");
        end

       1423 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1423");
        end

       1424 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1424");
        end

       1425 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1425");
        end

       1426 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1426");
        end

       1427 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1427");
        end

       1428 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1428");
        end

       1429 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1429");
        end

       1430 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1430");
        end

       1431 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1431");
        end

       1432 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1432");
        end

       1433 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1433");
        end

       1434 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1434");
        end

       1435 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1435");
        end

       1436 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1436");
        end

       1437 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1437");
        end

       1438 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1438");
        end

       1439 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1439");
        end

       1440 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1440");
        end

       1441 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1441");
        end

       1442 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1442");
        end

       1443 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1443");
        end

       1444 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1444");
        end

       1445 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1445");
        end

       1446 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1446");
        end

       1447 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1447");
        end

       1448 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1448");
        end

       1449 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1449");
        end

       1450 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1450");
        end

       1451 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1451");
        end

       1452 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1452");
        end

       1453 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1453");
        end

       1454 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1454");
        end

       1455 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1455");
        end

       1456 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1456");
        end

       1457 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1457");
        end

       1458 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1458");
        end

       1459 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1459");
        end

       1460 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1460");
        end

       1461 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1461");
        end

       1462 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1462");
        end

       1463 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1463");
        end

       1464 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1464");
        end

       1465 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1465");
        end

       1466 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1466");
        end

       1467 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1467");
        end

       1468 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1468");
        end

       1469 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1469");
        end

       1470 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1470");
        end

       1471 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1471");
        end

       1472 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1472");
        end

       1473 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1473");
        end

       1474 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1474");
        end

       1475 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1475");
        end

       1476 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1476");
        end

       1477 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1477");
        end

       1478 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1478");
        end

       1479 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1479");
        end

       1480 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1480");
        end

       1481 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1481");
        end

       1482 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1482");
        end

       1483 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1483");
        end

       1484 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1484");
        end

       1485 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1485");
        end

       1486 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1486");
        end

       1487 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1487");
        end

       1488 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1488");
        end

       1489 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1489");
        end

       1490 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1490");
        end

       1491 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1491");
        end

       1492 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1492");
        end

       1493 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1493");
        end

       1494 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1494");
        end

       1495 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1495");
        end

       1496 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1496");
        end

       1497 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1497");
        end

       1498 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1498");
        end

       1499 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1499");
        end

       1500 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1500");
        end

       1501 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1501");
        end

       1502 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1502");
        end

       1503 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1503");
        end

       1504 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1504");
        end

       1505 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1505");
        end

       1506 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1506");
        end

       1507 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1507");
        end

       1508 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1508");
        end

       1509 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1509");
        end

       1510 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1510");
        end

       1511 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1511");
        end

       1512 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1512");
        end

       1513 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1513");
        end

       1514 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1514");
        end

       1515 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1515");
        end

       1516 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1516");
        end

       1517 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1517");
        end

       1518 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1518");
        end

       1519 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1519");
        end

       1520 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1520");
        end

       1521 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1521");
        end

       1522 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1522");
        end

       1523 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1523");
        end

       1524 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1524");
        end

       1525 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1525");
        end

       1526 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1526");
        end

       1527 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1527");
        end

       1528 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1528");
        end

       1529 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1529");
        end

       1530 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1530");
        end

       1531 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1531");
        end

       1532 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1532");
        end

       1533 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1533");
        end

       1534 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1534");
        end

       1535 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1535");
        end

       1536 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1536");
        end

       1537 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1537");
        end

       1538 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1538");
        end

       1539 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1539");
        end

       1540 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1540");
        end

       1541 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1541");
        end

       1542 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1542");
        end

       1543 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1543");
        end

       1544 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1544");
        end

       1545 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1545");
        end

       1546 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1546");
        end

       1547 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1547");
        end

       1548 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1548");
        end

       1549 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1549");
        end

       1550 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1550");
        end

       1551 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1551");
        end

       1552 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1552");
        end

       1553 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1553");
        end

       1554 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1554");
        end

       1555 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1555");
        end

       1556 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1556");
        end

       1557 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1557");
        end

       1558 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1558");
        end

       1559 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1559");
        end

       1560 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1560");
        end

       1561 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1561");
        end

       1562 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1562");
        end

       1563 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1563");
        end

       1564 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1564");
        end

       1565 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1565");
        end

       1566 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1566");
        end

       1567 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1567");
        end

       1568 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1568");
        end

       1569 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1569");
        end

       1570 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1570");
        end

       1571 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1571");
        end

       1572 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1572");
        end

       1573 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1573");
        end

       1574 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1574");
        end

       1575 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1575");
        end

       1576 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1576");
        end

       1577 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1577");
        end

       1578 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1578");
        end

       1579 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1579");
        end

       1580 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1580");
        end

       1581 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1581");
        end

       1582 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1582");
        end

       1583 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1583");
        end

       1584 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1584");
        end

       1585 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1585");
        end

       1586 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1586");
        end

       1587 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1587");
        end

       1588 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1588");
        end

       1589 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1589");
        end

       1590 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1590");
        end

       1591 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1591");
        end

       1592 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1592");
        end

       1593 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1593");
        end

       1594 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1594");
        end

       1595 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1595");
        end

       1596 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1596");
        end

       1597 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1597");
        end

       1598 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1598");
        end

       1599 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1599");
        end

       1600 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1600");
        end

       1601 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1601");
        end

       1602 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1602");
        end

       1603 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1603");
        end

       1604 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1604");
        end

       1605 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1605");
        end

       1606 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1606");
        end

       1607 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1607");
        end

       1608 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1608");
        end

       1609 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1609");
        end

       1610 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1610");
        end

       1611 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1611");
        end

       1612 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1612");
        end

       1613 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1613");
        end

       1614 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1614");
        end

       1615 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1615");
        end

       1616 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1616");
        end

       1617 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1617");
        end

       1618 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1618");
        end

       1619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1619");
        end

       1620 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1620");
        end

       1621 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1621");
        end

       1622 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1622");
        end

       1623 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1623");
        end

       1624 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1624");
        end

       1625 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1625");
        end

       1626 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1626");
        end

       1627 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1627");
        end

       1628 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1628");
        end

       1629 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1629");
        end

       1630 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1630");
        end

       1631 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1631");
        end

       1632 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1632");
        end

       1633 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1633");
        end

       1634 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1634");
        end

       1635 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1635");
        end

       1636 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1636");
        end

       1637 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1637");
        end

       1638 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1638");
        end

       1639 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1639");
        end

       1640 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1640");
        end

       1641 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1641");
        end

       1642 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1642");
        end

       1643 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1643");
        end

       1644 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1644");
        end

       1645 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1645");
        end

       1646 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1646");
        end

       1647 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1647");
        end

       1648 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1648");
        end

       1649 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1649");
        end

       1650 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1650");
        end

       1651 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1651");
        end

       1652 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1652");
        end

       1653 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1653");
        end

       1654 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1654");
        end

       1655 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1655");
        end

       1656 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1656");
        end

       1657 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1657");
        end

       1658 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1658");
        end

       1659 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1659");
        end

       1660 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1660");
        end

       1661 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1661");
        end

       1662 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1662");
        end

       1663 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1663");
        end

       1664 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1664");
        end

       1665 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1665");
        end

       1666 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1666");
        end

       1667 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1667");
        end

       1668 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1668");
        end

       1669 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1669");
        end

       1670 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1670");
        end

       1671 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1671");
        end

       1672 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1672");
        end

       1673 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1673");
        end

       1674 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1674");
        end

       1675 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1675");
        end

       1676 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1676");
        end

       1677 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1677");
        end

       1678 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1678");
        end

       1679 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1679");
        end

       1680 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1680");
        end

       1681 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1681");
        end

       1682 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1682");
        end

       1683 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1683");
        end

       1684 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1684");
        end

       1685 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1686;
        end

       1686 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[142] = 1;
              ip = 1687;
        end

       1687 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1690;
        end

       1688 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1689;
        end

       1689 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[142] = 0;
              ip = 1690;
        end

       1690 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1691;
        end

       1691 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[142] != 0 ? 1693 : 1692;
        end

       1692 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[26] = localMem[141];
              ip = 1693;
        end

       1693 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1694;
        end

       1694 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2453;
        end

       1695 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1695");
        end

       1696 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1696");
        end

       1697 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1697");
        end

       1698 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1698");
        end

       1699 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1699");
        end

       1700 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1700");
        end

       1701 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1701");
        end

       1702 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1702");
        end

       1703 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1703");
        end

       1704 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1704");
        end

       1705 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1705");
        end

       1706 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1706");
        end

       1707 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1707");
        end

       1708 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1708");
        end

       1709 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1709");
        end

       1710 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1710");
        end

       1711 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1711");
        end

       1712 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1712");
        end

       1713 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1713");
        end

       1714 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1714");
        end

       1715 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1715");
        end

       1716 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed  1716");
        end

       1717 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1717");
        end

       1718 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1718");
        end

       1719 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1719");
        end

       1720 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1720");
        end

       1721 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1721");
        end

       1722 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1722");
        end

       1723 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1723");
        end

       1724 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1724");
        end

       1725 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1725");
        end

       1726 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1726");
        end

       1727 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1727");
        end

       1728 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1728");
        end

       1729 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1729");
        end

       1730 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1730");
        end

       1731 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1731");
        end

       1732 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1732");
        end

       1733 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1733");
        end

       1734 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1734");
        end

       1735 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1735");
        end

       1736 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1736");
        end

       1737 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1737");
        end

       1738 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1738");
        end

       1739 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1739");
        end

       1740 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1740");
        end

       1741 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1741");
        end

       1742 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1742");
        end

       1743 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1743");
        end

       1744 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1744");
        end

       1745 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1745");
        end

       1746 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1746");
        end

       1747 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1747");
        end

       1748 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1748");
        end

       1749 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1749");
        end

       1750 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1750");
        end

       1751 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1751");
        end

       1752 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1752");
        end

       1753 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1753");
        end

       1754 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1754");
        end

       1755 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1755");
        end

       1756 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1756");
        end

       1757 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1757");
        end

       1758 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1758");
        end

       1759 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1759");
        end

       1760 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1760");
        end

       1761 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1761");
        end

       1762 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
          // $display("Should not be executed  1762");
        end

       1763 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1763");
        end

       1764 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
          // $display("Should not be executed  1764");
        end

       1765 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1765");
        end

       1766 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1766");
        end

       1767 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1767");
        end

       1768 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1768");
        end

       1769 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1769");
        end

       1770 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1770");
        end

       1771 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1771");
        end

       1772 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1772");
        end

       1773 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1773");
        end

       1774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1774");
        end

       1775 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1775");
        end

       1776 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1776");
        end

       1777 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1777");
        end

       1778 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1778");
        end

       1779 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1779");
        end

       1780 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1780");
        end

       1781 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1781");
        end

       1782 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1782");
        end

       1783 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1783");
        end

       1784 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1784");
        end

       1785 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1785");
        end

       1786 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1786");
        end

       1787 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1787");
        end

       1788 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1788");
        end

       1789 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1789");
        end

       1790 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1790");
        end

       1791 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1791");
        end

       1792 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1792");
        end

       1793 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1793");
        end

       1794 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1794");
        end

       1795 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1795");
        end

       1796 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1796");
        end

       1797 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1797");
        end

       1798 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1798");
        end

       1799 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1799");
        end

       1800 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1800");
        end

       1801 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1801");
        end

       1802 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1802");
        end

       1803 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1803");
        end

       1804 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1804");
        end

       1805 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1805");
        end

       1806 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1806");
        end

       1807 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1807");
        end

       1808 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1808");
        end

       1809 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1809");
        end

       1810 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1810");
        end

       1811 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1811");
        end

       1812 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1812");
        end

       1813 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1813");
        end

       1814 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1814");
        end

       1815 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1815");
        end

       1816 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1816");
        end

       1817 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1817");
        end

       1818 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1818");
        end

       1819 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1819");
        end

       1820 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1820");
        end

       1821 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1821");
        end

       1822 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1822");
        end

       1823 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1823");
        end

       1824 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1824");
        end

       1825 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1825");
        end

       1826 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1826");
        end

       1827 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1827");
        end

       1828 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1828");
        end

       1829 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1829");
        end

       1830 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1830");
        end

       1831 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1831");
        end

       1832 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1832");
        end

       1833 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1833");
        end

       1834 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1834");
        end

       1835 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1835");
        end

       1836 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1836");
        end

       1837 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1837");
        end

       1838 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1838");
        end

       1839 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1839");
        end

       1840 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1840");
        end

       1841 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1841");
        end

       1842 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1842");
        end

       1843 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1843");
        end

       1844 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1844");
        end

       1845 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1845");
        end

       1846 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1846");
        end

       1847 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1847");
        end

       1848 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1848");
        end

       1849 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1849");
        end

       1850 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1850");
        end

       1851 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1851");
        end

       1852 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1852");
        end

       1853 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1853");
        end

       1854 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1854");
        end

       1855 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1855");
        end

       1856 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1856");
        end

       1857 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1857");
        end

       1858 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1858");
        end

       1859 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1859");
        end

       1860 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1860");
        end

       1861 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1861");
        end

       1862 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1862");
        end

       1863 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1863");
        end

       1864 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1864");
        end

       1865 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1865");
        end

       1866 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1866");
        end

       1867 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1867");
        end

       1868 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1868");
        end

       1869 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1869");
        end

       1870 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1870");
        end

       1871 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1871");
        end

       1872 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1872");
        end

       1873 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1873");
        end

       1874 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1874");
        end

       1875 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1875");
        end

       1876 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1876");
        end

       1877 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1877");
        end

       1878 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1878");
        end

       1879 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1879");
        end

       1880 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1880");
        end

       1881 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1881");
        end

       1882 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1882");
        end

       1883 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1883");
        end

       1884 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1884");
        end

       1885 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1885");
        end

       1886 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1886");
        end

       1887 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1887");
        end

       1888 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1888");
        end

       1889 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1889");
        end

       1890 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1890");
        end

       1891 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1891");
        end

       1892 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1892");
        end

       1893 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1893");
        end

       1894 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1894");
        end

       1895 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1895");
        end

       1896 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1896");
        end

       1897 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1897");
        end

       1898 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1898");
        end

       1899 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1899");
        end

       1900 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1900");
        end

       1901 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1901");
        end

       1902 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1902");
        end

       1903 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1903");
        end

       1904 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1904");
        end

       1905 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1905");
        end

       1906 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1906");
        end

       1907 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1907");
        end

       1908 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1908");
        end

       1909 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1909");
        end

       1910 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1910");
        end

       1911 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1911");
        end

       1912 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1912");
        end

       1913 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1913");
        end

       1914 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1914");
        end

       1915 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1915");
        end

       1916 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1916");
        end

       1917 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1917");
        end

       1918 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1918");
        end

       1919 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1919");
        end

       1920 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1920");
        end

       1921 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1921");
        end

       1922 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1922");
        end

       1923 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1923");
        end

       1924 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1924");
        end

       1925 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1925");
        end

       1926 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1926");
        end

       1927 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1927");
        end

       1928 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1928");
        end

       1929 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1929");
        end

       1930 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1930");
        end

       1931 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1931");
        end

       1932 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1932");
        end

       1933 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1933");
        end

       1934 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1934");
        end

       1935 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1935");
        end

       1936 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1936");
        end

       1937 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1937");
        end

       1938 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1938");
        end

       1939 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1939");
        end

       1940 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1940");
        end

       1941 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1941");
        end

       1942 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1942");
        end

       1943 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1943");
        end

       1944 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1944");
        end

       1945 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1945");
        end

       1946 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1946");
        end

       1947 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1947");
        end

       1948 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1948");
        end

       1949 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1949");
        end

       1950 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1950");
        end

       1951 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1951");
        end

       1952 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1952");
        end

       1953 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1953");
        end

       1954 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1954");
        end

       1955 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1955");
        end

       1956 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1956");
        end

       1957 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1957");
        end

       1958 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1958");
        end

       1959 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1959");
        end

       1960 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1960");
        end

       1961 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1961");
        end

       1962 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1962");
        end

       1963 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1963");
        end

       1964 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1964");
        end

       1965 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1965");
        end

       1966 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1966");
        end

       1967 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1967");
        end

       1968 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1968");
        end

       1969 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1969");
        end

       1970 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1970");
        end

       1971 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1971");
        end

       1972 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1972");
        end

       1973 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1973");
        end

       1974 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1974");
        end

       1975 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1975");
        end

       1976 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1976");
        end

       1977 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1977");
        end

       1978 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1978");
        end

       1979 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1979");
        end

       1980 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1980");
        end

       1981 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1981");
        end

       1982 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1982");
        end

       1983 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1983");
        end

       1984 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1984");
        end

       1985 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1985");
        end

       1986 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1986");
        end

       1987 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1987");
        end

       1988 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1988");
        end

       1989 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1989");
        end

       1990 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1990");
        end

       1991 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1991");
        end

       1992 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1992");
        end

       1993 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1993");
        end

       1994 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1994");
        end

       1995 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1995");
        end

       1996 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1996");
        end

       1997 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1997");
        end

       1998 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1998");
        end

       1999 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  1999");
        end

       2000 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2000");
        end

       2001 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2001");
        end

       2002 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2002");
        end

       2003 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2003");
        end

       2004 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2004");
        end

       2005 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2005");
        end

       2006 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2006");
        end

       2007 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  2007");
        end

       2008 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2008");
        end

       2009 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2009");
        end

       2010 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2010");
        end

       2011 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2011");
        end

       2012 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2012");
        end

       2013 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  2013");
        end

       2014 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2014");
        end

       2015 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2015");
        end

       2016 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  2016");
        end

       2017 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2017");
        end

       2018 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2018");
        end

       2019 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2019");
        end

       2020 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2020");
        end

       2021 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2021");
        end

       2022 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2022");
        end

       2023 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2023");
        end

       2024 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2024");
        end

       2025 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2025");
        end

       2026 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2026");
        end

       2027 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2027");
        end

       2028 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2028");
        end

       2029 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2029");
        end

       2030 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2030");
        end

       2031 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2031");
        end

       2032 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2032");
        end

       2033 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2033");
        end

       2034 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2034");
        end

       2035 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2035");
        end

       2036 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2036");
        end

       2037 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2037");
        end

       2038 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2038");
        end

       2039 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2039");
        end

       2040 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2040");
        end

       2041 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2041");
        end

       2042 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2042");
        end

       2043 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2043");
        end

       2044 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2044");
        end

       2045 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2045");
        end

       2046 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2046");
        end

       2047 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2047");
        end

       2048 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2048");
        end

       2049 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2049");
        end

       2050 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2050");
        end

       2051 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2051");
        end

       2052 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2052");
        end

       2053 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2053");
        end

       2054 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2054");
        end

       2055 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2055");
        end

       2056 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2056");
        end

       2057 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2057");
        end

       2058 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2058");
        end

       2059 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2059");
        end

       2060 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2060");
        end

       2061 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2061");
        end

       2062 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2062");
        end

       2063 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2063");
        end

       2064 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2064");
        end

       2065 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2065");
        end

       2066 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2066");
        end

       2067 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2067");
        end

       2068 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2068");
        end

       2069 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2069");
        end

       2070 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2070");
        end

       2071 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2071");
        end

       2072 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2072");
        end

       2073 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2073");
        end

       2074 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2074");
        end

       2075 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2075");
        end

       2076 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2076");
        end

       2077 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2077");
        end

       2078 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2078");
        end

       2079 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2079");
        end

       2080 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2080");
        end

       2081 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2081");
        end

       2082 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2082");
        end

       2083 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2083");
        end

       2084 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2084");
        end

       2085 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2085");
        end

       2086 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2086");
        end

       2087 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2087");
        end

       2088 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2088");
        end

       2089 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2089");
        end

       2090 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2090");
        end

       2091 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2091");
        end

       2092 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2092");
        end

       2093 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2093");
        end

       2094 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2094");
        end

       2095 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2095");
        end

       2096 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2096");
        end

       2097 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2097");
        end

       2098 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2098");
        end

       2099 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2099");
        end

       2100 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2100");
        end

       2101 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2101");
        end

       2102 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2102");
        end

       2103 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2103");
        end

       2104 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2104");
        end

       2105 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2105");
        end

       2106 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2106");
        end

       2107 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2107");
        end

       2108 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2108");
        end

       2109 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2109");
        end

       2110 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2110");
        end

       2111 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2111");
        end

       2112 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2112");
        end

       2113 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2113");
        end

       2114 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2114");
        end

       2115 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2115");
        end

       2116 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2116");
        end

       2117 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2117");
        end

       2118 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2118");
        end

       2119 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2119");
        end

       2120 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2120");
        end

       2121 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2121");
        end

       2122 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2122");
        end

       2123 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2123");
        end

       2124 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2124");
        end

       2125 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2125");
        end

       2126 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2126");
        end

       2127 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2127");
        end

       2128 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2128");
        end

       2129 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2129");
        end

       2130 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2130");
        end

       2131 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2131");
        end

       2132 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2132");
        end

       2133 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2133");
        end

       2134 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2134");
        end

       2135 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2135");
        end

       2136 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2136");
        end

       2137 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2137");
        end

       2138 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2138");
        end

       2139 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2139");
        end

       2140 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2140");
        end

       2141 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2141");
        end

       2142 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2142");
        end

       2143 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2143");
        end

       2144 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2144");
        end

       2145 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2145");
        end

       2146 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2146");
        end

       2147 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2147");
        end

       2148 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2148");
        end

       2149 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2149");
        end

       2150 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2150");
        end

       2151 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2151");
        end

       2152 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2152");
        end

       2153 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2153");
        end

       2154 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2154");
        end

       2155 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2155");
        end

       2156 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2156");
        end

       2157 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2157");
        end

       2158 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2158");
        end

       2159 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2159");
        end

       2160 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2160");
        end

       2161 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2161");
        end

       2162 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2162");
        end

       2163 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2163");
        end

       2164 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  2164");
        end

       2165 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  2165");
        end

       2166 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2166");
        end

       2167 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2167");
        end

       2168 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2168");
        end

       2169 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2169");
        end

       2170 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2170");
        end

       2171 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2171");
        end

       2172 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2172");
        end

       2173 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2173");
        end

       2174 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2174");
        end

       2175 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2175");
        end

       2176 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2176");
        end

       2177 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2177");
        end

       2178 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2178");
        end

       2179 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2179");
        end

       2180 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2180");
        end

       2181 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2181");
        end

       2182 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2182");
        end

       2183 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2183");
        end

       2184 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2184");
        end

       2185 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2185");
        end

       2186 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2186");
        end

       2187 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2187");
        end

       2188 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2188");
        end

       2189 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2189");
        end

       2190 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2190");
        end

       2191 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2191");
        end

       2192 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2192");
        end

       2193 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2193");
        end

       2194 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2194");
        end

       2195 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2195");
        end

       2196 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2196");
        end

       2197 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2197");
        end

       2198 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2198");
        end

       2199 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2199");
        end

       2200 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2200");
        end

       2201 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2201");
        end

       2202 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2202");
        end

       2203 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2203");
        end

       2204 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2204");
        end

       2205 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2205");
        end

       2206 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2206");
        end

       2207 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2207");
        end

       2208 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2208");
        end

       2209 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2209");
        end

       2210 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2210");
        end

       2211 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2211");
        end

       2212 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2212");
        end

       2213 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2213");
        end

       2214 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2214");
        end

       2215 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2215");
        end

       2216 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2216");
        end

       2217 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2217");
        end

       2218 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2218");
        end

       2219 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2219");
        end

       2220 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2220");
        end

       2221 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2221");
        end

       2222 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2222");
        end

       2223 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2223");
        end

       2224 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2224");
        end

       2225 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2225");
        end

       2226 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2226");
        end

       2227 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2227");
        end

       2228 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2228");
        end

       2229 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2229");
        end

       2230 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2230");
        end

       2231 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2231");
        end

       2232 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2232");
        end

       2233 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2233");
        end

       2234 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2234");
        end

       2235 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2235");
        end

       2236 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2236");
        end

       2237 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2237");
        end

       2238 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2238");
        end

       2239 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2239");
        end

       2240 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2240");
        end

       2241 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2241");
        end

       2242 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2242");
        end

       2243 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2243");
        end

       2244 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2244");
        end

       2245 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2245");
        end

       2246 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2246");
        end

       2247 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2247");
        end

       2248 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2248");
        end

       2249 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2249");
        end

       2250 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2250");
        end

       2251 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2251");
        end

       2252 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2252");
        end

       2253 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2253");
        end

       2254 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2254");
        end

       2255 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2255");
        end

       2256 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2256");
        end

       2257 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2257");
        end

       2258 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2258");
        end

       2259 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2259");
        end

       2260 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2260");
        end

       2261 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2261");
        end

       2262 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2262");
        end

       2263 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2263");
        end

       2264 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2264");
        end

       2265 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2265");
        end

       2266 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2266");
        end

       2267 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2267");
        end

       2268 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2268");
        end

       2269 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2269");
        end

       2270 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2270");
        end

       2271 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2271");
        end

       2272 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2272");
        end

       2273 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2273");
        end

       2274 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2274");
        end

       2275 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2275");
        end

       2276 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2276");
        end

       2277 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2277");
        end

       2278 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2278");
        end

       2279 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2279");
        end

       2280 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2280");
        end

       2281 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2281");
        end

       2282 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2282");
        end

       2283 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2283");
        end

       2284 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2284");
        end

       2285 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2285");
        end

       2286 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2286");
        end

       2287 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2287");
        end

       2288 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2288");
        end

       2289 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2289");
        end

       2290 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2290");
        end

       2291 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2291");
        end

       2292 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2292");
        end

       2293 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2293");
        end

       2294 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2294");
        end

       2295 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2295");
        end

       2296 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2296");
        end

       2297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2297");
        end

       2298 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2298");
        end

       2299 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2299");
        end

       2300 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2300");
        end

       2301 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2301");
        end

       2302 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2302");
        end

       2303 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2303");
        end

       2304 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2304");
        end

       2305 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2305");
        end

       2306 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2306");
        end

       2307 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2307");
        end

       2308 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2308");
        end

       2309 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2309");
        end

       2310 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2310");
        end

       2311 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2311");
        end

       2312 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2312");
        end

       2313 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2313");
        end

       2314 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2314");
        end

       2315 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2315");
        end

       2316 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2316");
        end

       2317 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2317");
        end

       2318 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2318");
        end

       2319 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2319");
        end

       2320 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2320");
        end

       2321 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2321");
        end

       2322 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2322");
        end

       2323 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2323");
        end

       2324 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2324");
        end

       2325 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2325");
        end

       2326 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2326");
        end

       2327 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2327");
        end

       2328 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2328");
        end

       2329 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2329");
        end

       2330 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2330");
        end

       2331 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2331");
        end

       2332 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2332");
        end

       2333 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2333");
        end

       2334 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2334");
        end

       2335 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2335");
        end

       2336 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2336");
        end

       2337 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2337");
        end

       2338 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2338");
        end

       2339 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2339");
        end

       2340 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2340");
        end

       2341 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2341");
        end

       2342 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2342");
        end

       2343 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2343");
        end

       2344 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2344");
        end

       2345 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2345");
        end

       2346 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2346");
        end

       2347 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2347");
        end

       2348 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2348");
        end

       2349 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2349");
        end

       2350 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2350");
        end

       2351 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2351");
        end

       2352 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2352");
        end

       2353 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2353");
        end

       2354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2354");
        end

       2355 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2355");
        end

       2356 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2356");
        end

       2357 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2357");
        end

       2358 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2358");
        end

       2359 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2359");
        end

       2360 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2360");
        end

       2361 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2361");
        end

       2362 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2362");
        end

       2363 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2363");
        end

       2364 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2364");
        end

       2365 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2365");
        end

       2366 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2366");
        end

       2367 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2367");
        end

       2368 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2368");
        end

       2369 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2369");
        end

       2370 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2370");
        end

       2371 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2371");
        end

       2372 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2372");
        end

       2373 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2373");
        end

       2374 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2374");
        end

       2375 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2375");
        end

       2376 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2376");
        end

       2377 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2377");
        end

       2378 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2378");
        end

       2379 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2379");
        end

       2380 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2380");
        end

       2381 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2381");
        end

       2382 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2382");
        end

       2383 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2383");
        end

       2384 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2384");
        end

       2385 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2385");
        end

       2386 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2386");
        end

       2387 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2387");
        end

       2388 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2388");
        end

       2389 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2389");
        end

       2390 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2390");
        end

       2391 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2391");
        end

       2392 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2392");
        end

       2393 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2393");
        end

       2394 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2394");
        end

       2395 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2395");
        end

       2396 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2396");
        end

       2397 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2397");
        end

       2398 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2398");
        end

       2399 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2399");
        end

       2400 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2400");
        end

       2401 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2401");
        end

       2402 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2402");
        end

       2403 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2403");
        end

       2404 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2404");
        end

       2405 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2405");
        end

       2406 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2406");
        end

       2407 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2407");
        end

       2408 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2408");
        end

       2409 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2409");
        end

       2410 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2410");
        end

       2411 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2411");
        end

       2412 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2412");
        end

       2413 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2413");
        end

       2414 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2414");
        end

       2415 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2415");
        end

       2416 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2416");
        end

       2417 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2417");
        end

       2418 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2418");
        end

       2419 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2419");
        end

       2420 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2420");
        end

       2421 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2421");
        end

       2422 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2422");
        end

       2423 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2423");
        end

       2424 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2424");
        end

       2425 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2425");
        end

       2426 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2426");
        end

       2427 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2427");
        end

       2428 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2428");
        end

       2429 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2429");
        end

       2430 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2430");
        end

       2431 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2431");
        end

       2432 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2432");
        end

       2433 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2433");
        end

       2434 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2434");
        end

       2435 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2435");
        end

       2436 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2436");
        end

       2437 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2437");
        end

       2438 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2438");
        end

       2439 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2439");
        end

       2440 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2440");
        end

       2441 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2441");
        end

       2442 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2442");
        end

       2443 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2443");
        end

       2444 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2444");
        end

       2445 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2445");
        end

       2446 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2446");
        end

       2447 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2447");
        end

       2448 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2448");
        end

       2449 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2449");
        end

       2450 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  2450");
        end

       2451 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2451");
        end

       2452 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2452");
        end

       2453 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2454;
        end

       2454 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[134] = localMem[134] + 1;
              ip = 2455;
        end

       2455 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 941;
        end

       2456 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2456");
        end

       2457 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  2457");
        end

       2458 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2458");
        end

       2459 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2459");
        end

       2460 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2461;
        end

       2461 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2462;
              heapClock = 1;
        end

       2462 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2463;
        end

       2463 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[970] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2464;
              heapClock = 1;
        end

       2464 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2465;
        end

       2465 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[362] = localMem[970];
              ip = 2466;
        end

       2466 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2467;
              heapClock = 1;
        end

       2467 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2468;
        end

       2468 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[971] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2469;
              heapClock = 1;
        end

       2469 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2470;
        end

       2470 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[363] = localMem[971];
              ip = 2471;
        end

       2471 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2472;
              heapClock = 1;
        end

       2472 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2473;
        end

       2473 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[972] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2474;
              heapClock = 1;
        end

       2474 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2475;
        end

       2475 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[364] = localMem[972];
              ip = 2476;
        end

       2476 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[363] != 1 ? 2486 : 2477;
        end

       2477 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2477");
        end

       2478 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2478");
        end

       2479 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2479");
        end

       2480 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2480");
        end

       2481 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2481");
        end

       2482 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2482");
        end

       2483 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2483");
        end

       2484 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2484");
        end

       2485 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2485");
        end

       2486 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2487;
        end

       2487 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[363] != 2 ? 2509 : 2488;
        end

       2488 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[366] = localMem[364] + 1;
              ip = 2489;
        end

       2489 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2490;
              heapClock = 1;
        end

       2490 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2491;
        end

       2491 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[975] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2492;
              heapClock = 1;
        end

       2492 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2493;
        end

       2493 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[367] = localMem[975];
              ip = 2494;
        end

       2494 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[1];
              heapArray  = localMem[367];
              heapIndex  = localMem[366];
              ip = 2495;
              heapClock = 1;
        end

       2495 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2496;
              heapClock = 1;
        end

       2496 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2497;
        end

       2497 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[976] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2498;
              heapClock = 1;
        end

       2498 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2499;
        end

       2499 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[368] = localMem[976];
              ip = 2500;
        end

       2500 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[2];
              heapArray  = localMem[368];
              heapIndex  = localMem[366];
              ip = 2501;
              heapClock = 1;
        end

       2501 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2502;
              heapClock = 1;
        end

       2502 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2503;
        end

       2503 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[977] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2504;
              heapClock = 1;
        end

       2504 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2505;
        end

       2505 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[978] = localMem[977] + 1;
              ip = 2506;
        end

       2506 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[362];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[978];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2507;
              heapClock = 1;
        end

       2507 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2508;
        end

       2508 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2529;
        end

       2509 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2509");
        end

       2510 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2510");
        end

       2511 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2511");
        end

       2512 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2512");
        end

       2513 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2513");
        end

       2514 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2514");
        end

       2515 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2515");
        end

       2516 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2516");
        end

       2517 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2517");
        end

       2518 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2518");
        end

       2519 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2519");
        end

       2520 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2520");
        end

       2521 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2521");
        end

       2522 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2522");
        end

       2523 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2523");
        end

       2524 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2524");
        end

       2525 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2525");
        end

       2526 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2526");
        end

       2527 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2527");
        end

       2528 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2528");
        end

       2529 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2530;
        end

       2530 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2531;
              heapClock = 1;
        end

       2531 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2532;
        end

       2532 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[983] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2533;
              heapClock = 1;
        end

       2533 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2534;
        end

       2534 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[984] = localMem[983] + 1;
              ip = 2535;
        end

       2535 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[984];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2536;
              heapClock = 1;
        end

       2536 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2537;
        end

       2537 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2538;
        end

       2538 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2539;
              heapClock = 1;
        end

       2539 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2540;
        end

       2540 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[985] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2541;
              heapClock = 1;
        end

       2541 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2542;
        end

       2542 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[372] = localMem[985];
              ip = 2543;
        end

       2543 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2544;
              heapClock = 1;
        end

       2544 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2545;
        end

       2545 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[986] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2546;
              heapClock = 1;
        end

       2546 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2547;
        end

       2547 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[373] = localMem[986];
              ip = 2548;
        end

       2548 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2549;
              heapClock = 1;
        end

       2549 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2550;
        end

       2550 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[987] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2551;
              heapClock = 1;
        end

       2551 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2552;
        end

       2552 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[374] = localMem[987];
              ip = 2553;
        end

       2553 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[372] <  localMem[374] ? 3238 : 2554;
        end

       2554 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[375] = localMem[374];
              ip = 2555;
        end

       2555 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
              localMem[375] = localMem[375] >> 1;
              ip = 2556;
              ip = 2556;
        end

       2556 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[376] = localMem[375] + 1;
              ip = 2557;
        end

       2557 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2558;
              heapClock = 1;
        end

       2558 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2559;
        end

       2559 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[988] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2560;
              heapClock = 1;
        end

       2560 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2561;
        end

       2561 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[377] = localMem[988];
              ip = 2562;
        end

       2562 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[377] == 0 ? 2868 : 2563;
        end

       2563 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2564;
              heapClock = 1;
        end

       2564 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[378] = heapOut;
              ip = 2565;
        end

       2565 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2566;
        end

       2566 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[989] = localMem[375];
              ip = 2567;
        end

       2567 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[989];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2568;
              heapClock = 1;
        end

       2568 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2569;
        end

       2569 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[990] = 0;
              ip = 2570;
        end

       2570 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[990];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2571;
              heapClock = 1;
        end

       2571 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2572;
        end

       2572 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2573;
              heapClock = 1;
        end

       2573 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[379] = heapOut;
              ip = 2574;
        end

       2574 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2575;
        end

       2575 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[991] = localMem[379];
              ip = 2576;
        end

       2576 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[991];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2577;
              heapClock = 1;
        end

       2577 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2578;
        end

       2578 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2579;
              heapClock = 1;
        end

       2579 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[380] = heapOut;
              ip = 2580;
        end

       2580 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2581;
        end

       2581 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[992] = localMem[380];
              ip = 2582;
        end

       2582 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[992];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2583;
              heapClock = 1;
        end

       2583 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2584;
        end

       2584 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[993] = 0;
              ip = 2585;
        end

       2585 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[993];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2586;
              heapClock = 1;
        end

       2586 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2587;
        end

       2587 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[994] = localMem[373];
              ip = 2588;
        end

       2588 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[994];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2589;
              heapClock = 1;
        end

       2589 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2590;
        end

       2590 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2591;
              heapClock = 1;
        end

       2591 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2592;
        end

       2592 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[995] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2593;
              heapClock = 1;
        end

       2593 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2594;
        end

       2594 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[996] = localMem[995] + 1;
              ip = 2595;
        end

       2595 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[373];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[996];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2596;
              heapClock = 1;
        end

       2596 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2597;
        end

       2597 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[373];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2598;
              heapClock = 1;
        end

       2598 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2599;
        end

       2599 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[997] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2600;
              heapClock = 1;
        end

       2600 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2601;
        end

       2601 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[998] = localMem[997];
              ip = 2602;
        end

       2602 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[998];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2603;
              heapClock = 1;
        end

       2603 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2604;
        end

       2604 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2605;
              heapClock = 1;
        end

       2605 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2606;
        end

       2606 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[999] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2607;
              heapClock = 1;
        end

       2607 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2608;
        end

       2608 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[381] = !localMem[999];
              ip = 2609;
        end

       2609 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[381] != 0 ? 2687 : 2610;
        end

       2610 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2610");
        end

       2611 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2611");
        end

       2612 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2612");
        end

       2613 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2613");
        end

       2614 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2614");
        end

       2615 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2615");
        end

       2616 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2616");
        end

       2617 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2617");
        end

       2618 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2618");
        end

       2619 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2619");
        end

       2620 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2620");
        end

       2621 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2621");
        end

       2622 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2622");
        end

       2623 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2623");
        end

       2624 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2624");
        end

       2625 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2625");
        end

       2626 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2626");
        end

       2627 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2627");
        end

       2628 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2628");
        end

       2629 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2629");
        end

       2630 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2630");
        end

       2631 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2631");
        end

       2632 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2632");
        end

       2633 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2633");
        end

       2634 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2634");
        end

       2635 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2635");
        end

       2636 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2636");
        end

       2637 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2637");
        end

       2638 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2638");
        end

       2639 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2639");
        end

       2640 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2640");
        end

       2641 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2641");
        end

       2642 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2642");
        end

       2643 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2643");
        end

       2644 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2644");
        end

       2645 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2645");
        end

       2646 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2646");
        end

       2647 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2647");
        end

       2648 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2648");
        end

       2649 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2649");
        end

       2650 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2650");
        end

       2651 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2651");
        end

       2652 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2652");
        end

       2653 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2653");
        end

       2654 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2654");
        end

       2655 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2655");
        end

       2656 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2656");
        end

       2657 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2657");
        end

       2658 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2658");
        end

       2659 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2659");
        end

       2660 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2660");
        end

       2661 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2661");
        end

       2662 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2662");
        end

       2663 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2663");
        end

       2664 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2664");
        end

       2665 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2665");
        end

       2666 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2666");
        end

       2667 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2667");
        end

       2668 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2668");
        end

       2669 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2669");
        end

       2670 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2670");
        end

       2671 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2671");
        end

       2672 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2672");
        end

       2673 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2673");
        end

       2674 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2674");
        end

       2675 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2675");
        end

       2676 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2676");
        end

       2677 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2677");
        end

       2678 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2678");
        end

       2679 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2679");
        end

       2680 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2680");
        end

       2681 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2681");
        end

       2682 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2682");
        end

       2683 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2683");
        end

       2684 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2684");
        end

       2685 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2685");
        end

       2686 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2686");
        end

       2687 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2688;
        end

       2688 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2689;
              heapClock = 1;
        end

       2689 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2690;
        end

       2690 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1012] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2691;
              heapClock = 1;
        end

       2691 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2692;
        end

       2692 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[396] = localMem[1012];
              ip = 2693;
        end

       2693 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[378];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2694;
              heapClock = 1;
        end

       2694 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2695;
        end

       2695 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1013] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2696;
              heapClock = 1;
        end

       2696 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2697;
        end

       2697 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[397] = localMem[1013];
              ip = 2698;
        end

       2698 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[396];                                                 // Array to write to
              heapIndex  = localMem[376];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 2699;
              heapClock = 1;
        end

       2699 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[397];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[375];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 2700;
              heapClock = 1;
        end

       2700 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2701;
              heapClock = 1;
        end

       2701 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2702;
        end

       2702 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1014] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2703;
              heapClock = 1;
        end

       2703 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2704;
        end

       2704 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[398] = localMem[1014];
              ip = 2705;
        end

       2705 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[378];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2706;
              heapClock = 1;
        end

       2706 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2707;
        end

       2707 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1015] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2708;
              heapClock = 1;
        end

       2708 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2709;
        end

       2709 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[399] = localMem[1015];
              ip = 2710;
        end

       2710 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[398];                                                 // Array to write to
              heapIndex  = localMem[376];                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 2711;
              heapClock = 1;
        end

       2711 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[399];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[375];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 2712;
              heapClock = 1;
        end

       2712 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2713;
        end

       2713 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1016] = localMem[375];
              ip = 2714;
        end

       2714 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[362];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1016];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2715;
              heapClock = 1;
        end

       2715 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2716;
        end

       2716 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1017] = localMem[377];
              ip = 2717;
        end

       2717 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[378];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1017];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2718;
              heapClock = 1;
        end

       2718 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2719;
        end

       2719 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2720;
              heapClock = 1;
        end

       2720 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2721;
        end

       2721 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1018] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2722;
              heapClock = 1;
        end

       2722 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2723;
        end

       2723 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[400] = localMem[1018];
              ip = 2724;
        end

       2724 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2725;
              heapClock = 1;
        end

       2725 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2726;
        end

       2726 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1019] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2727;
              heapClock = 1;
        end

       2727 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2728;
        end

       2728 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[401] = localMem[1019];
              ip = 2729;
        end

       2729 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[401];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[400];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2730;
              heapClock = 1;
        end

       2730 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2731;
        end

       2731 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1020] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2732;
              heapClock = 1;
        end

       2732 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2733;
        end

       2733 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[402] = localMem[1020];
              ip = 2734;
        end

       2734 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[402] != localMem[362] ? 2797 : 2735;
        end

       2735 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2736;
              heapClock = 1;
        end

       2736 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2737;
        end

       2737 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1021] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2738;
              heapClock = 1;
        end

       2738 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2739;
        end

       2739 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[403] = localMem[1021];
              ip = 2740;
        end

       2740 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[403];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[375];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2741;
              heapClock = 1;
        end

       2741 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2742;
        end

       2742 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1022] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2743;
              heapClock = 1;
        end

       2743 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2744;
        end

       2744 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[404] = localMem[1022];
              ip = 2745;
        end

       2745 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2746;
              heapClock = 1;
        end

       2746 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2747;
        end

       2747 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1023] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2748;
              heapClock = 1;
        end

       2748 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2749;
        end

       2749 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[405] = localMem[1023];
              ip = 2750;
        end

       2750 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1024] = localMem[404];
              ip = 2751;
        end

       2751 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[405];                                                // Array to write to
              heapIndex   = localMem[400];                                                // Index of element to write to
              heapIn      = localMem[1024];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2752;
              heapClock = 1;
        end

       2752 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2753;
        end

       2753 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2754;
              heapClock = 1;
        end

       2754 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2755;
        end

       2755 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1025] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2756;
              heapClock = 1;
        end

       2756 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2757;
        end

       2757 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[406] = localMem[1025];
              ip = 2758;
        end

       2758 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[406];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[375];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2759;
              heapClock = 1;
        end

       2759 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2760;
        end

       2760 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1026] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2761;
              heapClock = 1;
        end

       2761 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2762;
        end

       2762 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[407] = localMem[1026];
              ip = 2763;
        end

       2763 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2764;
              heapClock = 1;
        end

       2764 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2765;
        end

       2765 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1027] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2766;
              heapClock = 1;
        end

       2766 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2767;
        end

       2767 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[408] = localMem[1027];
              ip = 2768;
        end

       2768 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1028] = localMem[407];
              ip = 2769;
        end

       2769 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[408];                                                // Array to write to
              heapIndex   = localMem[400];                                                // Index of element to write to
              heapIn      = localMem[1028];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2770;
              heapClock = 1;
        end

       2770 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2771;
        end

       2771 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2772;
              heapClock = 1;
        end

       2772 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2773;
        end

       2773 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1029] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2774;
              heapClock = 1;
        end

       2774 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2775;
        end

       2775 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[409] = localMem[1029];
              ip = 2776;
        end

       2776 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[375];
              heapArray  = localMem[409];
              ip = 2777;
              heapClock = 1;
        end

       2777 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[362];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2778;
              heapClock = 1;
        end

       2778 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2779;
        end

       2779 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1030] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2780;
              heapClock = 1;
        end

       2780 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2781;
        end

       2781 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[410] = localMem[1030];
              ip = 2782;
        end

       2782 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[375];
              heapArray  = localMem[410];
              ip = 2783;
              heapClock = 1;
        end

       2783 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[411] = localMem[400] + 1;
              ip = 2784;
        end

       2784 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1031] = localMem[411];
              ip = 2785;
        end

       2785 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[377];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1031];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2786;
              heapClock = 1;
        end

       2786 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2787;
        end

       2787 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[377];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2788;
              heapClock = 1;
        end

       2788 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2789;
        end

       2789 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1032] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2790;
              heapClock = 1;
        end

       2790 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2791;
        end

       2791 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[412] = localMem[1032];
              ip = 2792;
        end

       2792 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1033] = localMem[378];
              ip = 2793;
        end

       2793 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[412];                                                // Array to write to
              heapIndex   = localMem[411];                                                // Index of element to write to
              heapIn      = localMem[1033];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2794;
              heapClock = 1;
        end

       2794 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 2795;
        end

       2795 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3235;
        end

       2796 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2796");
        end

       2797 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2797");
        end

       2798 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  2798");
        end

       2799 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2799");
        end

       2800 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2800");
        end

       2801 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2801");
        end

       2802 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2802");
        end

       2803 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2803");
        end

       2804 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  2804");
        end

       2805 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2805");
        end

       2806 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2806");
        end

       2807 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  2807");
        end

       2808 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2808");
        end

       2809 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2809");
        end

       2810 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2810");
        end

       2811 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2811");
        end

       2812 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2812");
        end

       2813 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2813");
        end

       2814 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2814");
        end

       2815 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2815");
        end

       2816 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2816");
        end

       2817 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2817");
        end

       2818 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2818");
        end

       2819 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2819");
        end

       2820 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2820");
        end

       2821 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2821");
        end

       2822 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2822");
        end

       2823 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2823");
        end

       2824 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2824");
        end

       2825 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2825");
        end

       2826 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2826");
        end

       2827 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2827");
        end

       2828 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2828");
        end

       2829 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2829");
        end

       2830 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2830");
        end

       2831 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2831");
        end

       2832 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2832");
        end

       2833 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2833");
        end

       2834 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2834");
        end

       2835 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2835");
        end

       2836 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2836");
        end

       2837 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2837");
        end

       2838 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2838");
        end

       2839 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2839");
        end

       2840 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2840");
        end

       2841 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2841");
        end

       2842 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2842");
        end

       2843 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2843");
        end

       2844 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2844");
        end

       2845 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2845");
        end

       2846 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2846");
        end

       2847 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2847");
        end

       2848 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2848");
        end

       2849 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2849");
        end

       2850 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2850");
        end

       2851 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2851");
        end

       2852 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2852");
        end

       2853 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2853");
        end

       2854 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2854");
        end

       2855 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2855");
        end

       2856 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2856");
        end

       2857 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2857");
        end

       2858 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  2858");
        end

       2859 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2859");
        end

       2860 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2860");
        end

       2861 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2861");
        end

       2862 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2862");
        end

       2863 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2863");
        end

       2864 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2864");
        end

       2865 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2865");
        end

       2866 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2866");
        end

       2867 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2867");
        end

       2868 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2868");
        end

       2869 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2869");
        end

       2870 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2870");
        end

       2871 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2871");
        end

       2872 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2872");
        end

       2873 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2873");
        end

       2874 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2874");
        end

       2875 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2875");
        end

       2876 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2876");
        end

       2877 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2877");
        end

       2878 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2878");
        end

       2879 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2879");
        end

       2880 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2880");
        end

       2881 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2881");
        end

       2882 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2882");
        end

       2883 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2883");
        end

       2884 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2884");
        end

       2885 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2885");
        end

       2886 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2886");
        end

       2887 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2887");
        end

       2888 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2888");
        end

       2889 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2889");
        end

       2890 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2890");
        end

       2891 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2891");
        end

       2892 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2892");
        end

       2893 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2893");
        end

       2894 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2894");
        end

       2895 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2895");
        end

       2896 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2896");
        end

       2897 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2897");
        end

       2898 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2898");
        end

       2899 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2899");
        end

       2900 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2900");
        end

       2901 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2901");
        end

       2902 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2902");
        end

       2903 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2903");
        end

       2904 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2904");
        end

       2905 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2905");
        end

       2906 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2906");
        end

       2907 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2907");
        end

       2908 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2908");
        end

       2909 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2909");
        end

       2910 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2910");
        end

       2911 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2911");
        end

       2912 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2912");
        end

       2913 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2913");
        end

       2914 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2914");
        end

       2915 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2915");
        end

       2916 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2916");
        end

       2917 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2917");
        end

       2918 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2918");
        end

       2919 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2919");
        end

       2920 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2920");
        end

       2921 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2921");
        end

       2922 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2922");
        end

       2923 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2923");
        end

       2924 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2924");
        end

       2925 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2925");
        end

       2926 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2926");
        end

       2927 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2927");
        end

       2928 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2928");
        end

       2929 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2929");
        end

       2930 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2930");
        end

       2931 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2931");
        end

       2932 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2932");
        end

       2933 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2933");
        end

       2934 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2934");
        end

       2935 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2935");
        end

       2936 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2936");
        end

       2937 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2937");
        end

       2938 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2938");
        end

       2939 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2939");
        end

       2940 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2940");
        end

       2941 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2941");
        end

       2942 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2942");
        end

       2943 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2943");
        end

       2944 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2944");
        end

       2945 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2945");
        end

       2946 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2946");
        end

       2947 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2947");
        end

       2948 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2948");
        end

       2949 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2949");
        end

       2950 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2950");
        end

       2951 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2951");
        end

       2952 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2952");
        end

       2953 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2953");
        end

       2954 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2954");
        end

       2955 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  2955");
        end

       2956 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  2956");
        end

       2957 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2957");
        end

       2958 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2958");
        end

       2959 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2959");
        end

       2960 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2960");
        end

       2961 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2961");
        end

       2962 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2962");
        end

       2963 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2963");
        end

       2964 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2964");
        end

       2965 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2965");
        end

       2966 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2966");
        end

       2967 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2967");
        end

       2968 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2968");
        end

       2969 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2969");
        end

       2970 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2970");
        end

       2971 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2971");
        end

       2972 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2972");
        end

       2973 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2973");
        end

       2974 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2974");
        end

       2975 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2975");
        end

       2976 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2976");
        end

       2977 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2977");
        end

       2978 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2978");
        end

       2979 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2979");
        end

       2980 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2980");
        end

       2981 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2981");
        end

       2982 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2982");
        end

       2983 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2983");
        end

       2984 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2984");
        end

       2985 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2985");
        end

       2986 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2986");
        end

       2987 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2987");
        end

       2988 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2988");
        end

       2989 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2989");
        end

       2990 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2990");
        end

       2991 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2991");
        end

       2992 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2992");
        end

       2993 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2993");
        end

       2994 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2994");
        end

       2995 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2995");
        end

       2996 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2996");
        end

       2997 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2997");
        end

       2998 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2998");
        end

       2999 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  2999");
        end

       3000 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3000");
        end

       3001 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3001");
        end

       3002 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3002");
        end

       3003 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3003");
        end

       3004 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3004");
        end

       3005 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3005");
        end

       3006 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3006");
        end

       3007 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3007");
        end

       3008 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3008");
        end

       3009 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3009");
        end

       3010 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3010");
        end

       3011 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3011");
        end

       3012 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3012");
        end

       3013 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3013");
        end

       3014 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3014");
        end

       3015 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3015");
        end

       3016 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3016");
        end

       3017 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3017");
        end

       3018 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3018");
        end

       3019 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3019");
        end

       3020 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3020");
        end

       3021 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3021");
        end

       3022 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3022");
        end

       3023 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3023");
        end

       3024 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3024");
        end

       3025 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3025");
        end

       3026 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3026");
        end

       3027 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3027");
        end

       3028 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3028");
        end

       3029 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3029");
        end

       3030 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3030");
        end

       3031 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3031");
        end

       3032 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3032");
        end

       3033 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3033");
        end

       3034 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3034");
        end

       3035 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3035");
        end

       3036 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3036");
        end

       3037 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3037");
        end

       3038 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3038");
        end

       3039 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3039");
        end

       3040 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3040");
        end

       3041 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3041");
        end

       3042 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3042");
        end

       3043 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3043");
        end

       3044 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3044");
        end

       3045 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3045");
        end

       3046 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3046");
        end

       3047 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3047");
        end

       3048 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3048");
        end

       3049 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3049");
        end

       3050 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3050");
        end

       3051 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3051");
        end

       3052 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3052");
        end

       3053 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3053");
        end

       3054 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3054");
        end

       3055 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3055");
        end

       3056 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3056");
        end

       3057 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  3057");
        end

       3058 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3058");
        end

       3059 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3059");
        end

       3060 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3060");
        end

       3061 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3061");
        end

       3062 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3062");
        end

       3063 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3063");
        end

       3064 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3064");
        end

       3065 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3065");
        end

       3066 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3066");
        end

       3067 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3067");
        end

       3068 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3068");
        end

       3069 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3069");
        end

       3070 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3070");
        end

       3071 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3071");
        end

       3072 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3072");
        end

       3073 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3073");
        end

       3074 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3074");
        end

       3075 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3075");
        end

       3076 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3076");
        end

       3077 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3077");
        end

       3078 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3078");
        end

       3079 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3079");
        end

       3080 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3080");
        end

       3081 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3081");
        end

       3082 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3082");
        end

       3083 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3083");
        end

       3084 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  3084");
        end

       3085 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3085");
        end

       3086 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3086");
        end

       3087 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3087");
        end

       3088 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3088");
        end

       3089 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3089");
        end

       3090 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3090");
        end

       3091 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3091");
        end

       3092 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3092");
        end

       3093 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3093");
        end

       3094 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  3094");
        end

       3095 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3095");
        end

       3096 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3096");
        end

       3097 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3097");
        end

       3098 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3098");
        end

       3099 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  3099");
        end

       3100 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3100");
        end

       3101 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3101");
        end

       3102 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3102");
        end

       3103 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3103");
        end

       3104 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3104");
        end

       3105 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3105");
        end

       3106 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3106");
        end

       3107 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3107");
        end

       3108 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3108");
        end

       3109 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3109");
        end

       3110 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3110");
        end

       3111 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3111");
        end

       3112 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3112");
        end

       3113 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3113");
        end

       3114 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3114");
        end

       3115 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3115");
        end

       3116 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3116");
        end

       3117 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3117");
        end

       3118 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3118");
        end

       3119 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3119");
        end

       3120 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3120");
        end

       3121 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3121");
        end

       3122 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3122");
        end

       3123 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3123");
        end

       3124 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3124");
        end

       3125 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3125");
        end

       3126 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3126");
        end

       3127 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3127");
        end

       3128 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3128");
        end

       3129 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3129");
        end

       3130 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3130");
        end

       3131 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3131");
        end

       3132 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3132");
        end

       3133 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3133");
        end

       3134 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3134");
        end

       3135 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3135");
        end

       3136 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3136");
        end

       3137 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3137");
        end

       3138 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3138");
        end

       3139 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3139");
        end

       3140 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3140");
        end

       3141 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3141");
        end

       3142 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3142");
        end

       3143 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3143");
        end

       3144 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3144");
        end

       3145 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3145");
        end

       3146 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3146");
        end

       3147 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3147");
        end

       3148 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3148");
        end

       3149 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3149");
        end

       3150 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3150");
        end

       3151 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  3151");
        end

       3152 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  3152");
        end

       3153 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3153");
        end

       3154 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3154");
        end

       3155 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3155");
        end

       3156 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3156");
        end

       3157 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3157");
        end

       3158 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3158");
        end

       3159 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3159");
        end

       3160 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3160");
        end

       3161 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3161");
        end

       3162 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3162");
        end

       3163 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3163");
        end

       3164 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3164");
        end

       3165 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3165");
        end

       3166 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3166");
        end

       3167 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3167");
        end

       3168 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3168");
        end

       3169 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3169");
        end

       3170 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3170");
        end

       3171 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3171");
        end

       3172 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3172");
        end

       3173 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3173");
        end

       3174 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3174");
        end

       3175 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3175");
        end

       3176 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3176");
        end

       3177 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3177");
        end

       3178 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3178");
        end

       3179 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3179");
        end

       3180 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3180");
        end

       3181 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3181");
        end

       3182 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3182");
        end

       3183 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3183");
        end

       3184 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3184");
        end

       3185 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3185");
        end

       3186 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3186");
        end

       3187 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3187");
        end

       3188 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3188");
        end

       3189 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3189");
        end

       3190 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3190");
        end

       3191 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3191");
        end

       3192 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3192");
        end

       3193 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3193");
        end

       3194 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3194");
        end

       3195 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3195");
        end

       3196 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3196");
        end

       3197 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3197");
        end

       3198 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3198");
        end

       3199 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3199");
        end

       3200 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3200");
        end

       3201 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3201");
        end

       3202 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3202");
        end

       3203 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3203");
        end

       3204 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3204");
        end

       3205 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3205");
        end

       3206 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3206");
        end

       3207 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3207");
        end

       3208 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3208");
        end

       3209 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3209");
        end

       3210 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3210");
        end

       3211 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3211");
        end

       3212 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3212");
        end

       3213 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3213");
        end

       3214 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3214");
        end

       3215 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3215");
        end

       3216 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3216");
        end

       3217 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3217");
        end

       3218 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3218");
        end

       3219 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3219");
        end

       3220 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3220");
        end

       3221 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3221");
        end

       3222 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3222");
        end

       3223 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3223");
        end

       3224 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3224");
        end

       3225 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3225");
        end

       3226 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3226");
        end

       3227 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3227");
        end

       3228 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3228");
        end

       3229 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3229");
        end

       3230 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3230");
        end

       3231 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3231");
        end

       3232 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  3232");
        end

       3233 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3233");
        end

       3234 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3234");
        end

       3235 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3236;
        end

       3236 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[371] = 1;
              ip = 3237;
        end

       3237 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3240;
        end

       3238 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3239;
        end

       3239 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[371] = 0;
              ip = 3240;
        end

       3240 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3241;
        end

       3241 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3242;
        end

       3242 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3243;
        end

       3243 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3244;
        end

       3244 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[3];
              ip = 3245;
              heapClock = 1;
        end

       3245 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3246;
        end

       3246 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1] = localMem[1] + 1;
              ip = 3247;
        end

       3247 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 20;
        end

       3248 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3249;
        end

       3249 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3250;
        end

       3250 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[478] = 0;
              ip = 3251;
        end

       3251 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3252;
        end

       3252 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[478] >= 66 ? 3402 : 3253;
        end

       3253 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3254;
              heapClock = 1;
        end

       3254 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[479] = heapOut;
              ip = 3255;
        end

       3255 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3256;
        end

       3256 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3257;
        end

       3257 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3258;
              heapClock = 1;
        end

       3258 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3259;
        end

       3259 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1116] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3260;
              heapClock = 1;
        end

       3260 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3261;
        end

       3261 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[480] = localMem[1116];
              ip = 3262;
        end

       3262 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[480] != 0 ? 3273 : 3263;
        end

       3263 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3263");
        end

       3264 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3264");
        end

       3265 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3265");
        end

       3266 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3266");
        end

       3267 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3267");
        end

       3268 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3268");
        end

       3269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3269");
        end

       3270 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3270");
        end

       3271 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3271");
        end

       3272 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3272");
        end

       3273 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3274;
        end

       3274 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3275;
        end

       3275 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = 0;
              ip = 3276;
        end

       3276 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3277;
        end

       3277 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[481] >= 99 ? 3373 : 3278;
        end

       3278 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3279;
              heapClock = 1;
        end

       3279 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3280;
        end

       3280 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1120] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3281;
              heapClock = 1;
        end

       3281 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3282;
        end

       3282 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[482] = localMem[1120] - 1;
              ip = 3283;
        end

       3283 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3284;
              heapClock = 1;
        end

       3284 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3285;
        end

       3285 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1121] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3286;
              heapClock = 1;
        end

       3286 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3287;
        end

       3287 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[483] = localMem[1121];
              ip = 3288;
        end

       3288 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[483];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[482];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3289;
              heapClock = 1;
        end

       3289 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3290;
        end

       3290 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1122] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3291;
              heapClock = 1;
        end

       3291 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3292;
        end

       3292 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[478] <= localMem[1122] ? 3323 : 3293;
        end

       3293 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[484] = localMem[482] + 1;
              ip = 3294;
        end

       3294 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3295;
              heapClock = 1;
        end

       3295 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3296;
        end

       3296 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1123] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3297;
              heapClock = 1;
        end

       3297 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3298;
        end

       3298 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[485] = !localMem[1123];
              ip = 3299;
        end

       3299 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[485] == 0 ? 3310 : 3300;
        end

       3300 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3300");
        end

       3301 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3301");
        end

       3302 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3302");
        end

       3303 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3303");
        end

       3304 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3304");
        end

       3305 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3305");
        end

       3306 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3306");
        end

       3307 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3307");
        end

       3308 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3308");
        end

       3309 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3309");
        end

       3310 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3311;
        end

       3311 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3312;
              heapClock = 1;
        end

       3312 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3313;
        end

       3313 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1127] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3314;
              heapClock = 1;
        end

       3314 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3315;
        end

       3315 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[486] = localMem[1127];
              ip = 3316;
        end

       3316 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[486];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[484];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3317;
              heapClock = 1;
        end

       3317 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3318;
        end

       3318 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1128] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3319;
              heapClock = 1;
        end

       3319 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3320;
        end

       3320 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[487] = localMem[1128];
              ip = 3321;
        end

       3321 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[480] = localMem[487];
              ip = 3322;
        end

       3322 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3370;
        end

       3323 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3324;
        end

       3324 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[478];
              heapAction = `Index;
              heapArray  = localMem[483];
              ip = 3325;
              heapClock = 1;
        end

       3325 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[488] = heapOut;
              ip = 3326;
        end

       3326 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3327;
        end

       3327 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[488] == 0 ? 3338 : 3328;
        end

       3328 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1129] = localMem[480];
              ip = 3329;
        end

       3329 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[479];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1129];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3330;
              heapClock = 1;
        end

       3330 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3331;
        end

       3331 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1130] = 1;
              ip = 3332;
        end

       3332 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[479];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1130];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3333;
              heapClock = 1;
        end

       3333 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3334;
        end

       3334 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[1131] = localMem[488] - 1;
              ip = 3335;
        end

       3335 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[479];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1131];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3336;
              heapClock = 1;
        end

       3336 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3337;
        end

       3337 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3377;
        end

       3338 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3339;
        end

       3339 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
              heapIn     = localMem[478];
              heapAction = `Less;
              heapArray  = localMem[483];
              ip = 3340;
              heapClock = 1;
        end

       3340 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[489] = heapOut;
              ip = 3341;
        end

       3341 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3342;
        end

       3342 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3343;
              heapClock = 1;
        end

       3343 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3344;
        end

       3344 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1132] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3345;
              heapClock = 1;
        end

       3345 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3346;
        end

       3346 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[490] = !localMem[1132];
              ip = 3347;
        end

       3347 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[490] == 0 ? 3358 : 3348;
        end

       3348 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3348");
        end

       3349 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3349");
        end

       3350 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3350");
        end

       3351 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3351");
        end

       3352 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3352");
        end

       3353 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3353");
        end

       3354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3354");
        end

       3355 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3355");
        end

       3356 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3356");
        end

       3357 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3357");
        end

       3358 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3359;
        end

       3359 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[480];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3360;
              heapClock = 1;
        end

       3360 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3361;
        end

       3361 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1136] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3362;
              heapClock = 1;
        end

       3362 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3363;
        end

       3363 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[491] = localMem[1136];
              ip = 3364;
        end

       3364 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[491];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[489];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3365;
              heapClock = 1;
        end

       3365 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3366;
        end

       3366 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1137] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3367;
              heapClock = 1;
        end

       3367 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3368;
        end

       3368 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[492] = localMem[1137];
              ip = 3369;
        end

       3369 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[480] = localMem[492];
              ip = 3370;
        end

       3370 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3371;
        end

       3371 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[481] = localMem[481] + 1;
              ip = 3372;
        end

       3372 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3276;
        end

       3373 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3373");
        end

       3374 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  3374");
        end

       3375 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3375");
        end

       3376 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3376");
        end

       3377 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3378;
        end

       3378 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[479];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3379;
              heapClock = 1;
        end

       3379 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3380;
        end

       3380 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1138] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3381;
              heapClock = 1;
        end

       3381 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3382;
        end

       3382 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[493] = localMem[1138];
              ip = 3383;
        end

       3383 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[479];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3384;
              heapClock = 1;
        end

       3384 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3385;
        end

       3385 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1139] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3386;
              heapClock = 1;
        end

       3386 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3387;
        end

       3387 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[494] = localMem[1139];
              ip = 3388;
        end

       3388 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[493];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3389;
              heapClock = 1;
        end

       3389 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3390;
        end

       3390 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1140] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3391;
              heapClock = 1;
        end

       3391 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3392;
        end

       3392 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[495] = localMem[1140];
              ip = 3393;
        end

       3393 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[495];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[494];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3394;
              heapClock = 1;
        end

       3394 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3395;
        end

       3395 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1141] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3396;
              heapClock = 1;
        end

       3396 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3397;
        end

       3397 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[496] = localMem[1141];
              ip = 3398;
        end

       3398 :
        begin                                                                   // out
          //$display("AAAA %4d %4d out", steps, ip);
              outMem[outMemPos] = localMem[496];
              outMemPos = outMemPos + 1;
              ip = 3399;
        end

       3399 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3400;
        end

       3400 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[478] = localMem[478] + 1;
              ip = 3401;
        end

       3401 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3251;
        end

       3402 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3403;
        end

       3403 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3404;
              heapClock = 1;
        end

       3404 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[497] = heapOut;
              ip = 3405;
        end

       3405 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3406;
        end

       3406 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3407;
        end

       3407 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3408;
              heapClock = 1;
        end

       3408 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3409;
        end

       3409 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1142] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3410;
              heapClock = 1;
        end

       3410 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3411;
        end

       3411 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[498] = localMem[1142];
              ip = 3412;
        end

       3412 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[498] != 0 ? 3423 : 3413;
        end

       3413 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3413");
        end

       3414 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3414");
        end

       3415 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3415");
        end

       3416 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3416");
        end

       3417 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3417");
        end

       3418 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3418");
        end

       3419 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3419");
        end

       3420 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3420");
        end

       3421 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3421");
        end

       3422 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3422");
        end

       3423 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3424;
        end

       3424 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3425;
        end

       3425 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[499] = 0;
              ip = 3426;
        end

       3426 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3427;
        end

       3427 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[499] >= 99 ? 3523 : 3428;
        end

       3428 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3429;
              heapClock = 1;
        end

       3429 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3430;
        end

       3430 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1146] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3431;
              heapClock = 1;
        end

       3431 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3432;
        end

       3432 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[500] = localMem[1146] - 1;
              ip = 3433;
        end

       3433 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3434;
              heapClock = 1;
        end

       3434 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3435;
        end

       3435 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1147] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3436;
              heapClock = 1;
        end

       3436 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3437;
        end

       3437 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[501] = localMem[1147];
              ip = 3438;
        end

       3438 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[501];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[500];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3439;
              heapClock = 1;
        end

       3439 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3440;
        end

       3440 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1148] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3441;
              heapClock = 1;
        end

       3441 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3442;
        end

       3442 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = 66 <= localMem[1148] ? 3473 : 3443;
        end

       3443 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[502] = localMem[500] + 1;
              ip = 3444;
        end

       3444 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3445;
              heapClock = 1;
        end

       3445 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3446;
        end

       3446 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1149] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3447;
              heapClock = 1;
        end

       3447 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3448;
        end

       3448 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[503] = !localMem[1149];
              ip = 3449;
        end

       3449 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[503] == 0 ? 3460 : 3450;
        end

       3450 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1150] = localMem[498];
              ip = 3451;
        end

       3451 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[497];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1150];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3452;
              heapClock = 1;
        end

       3452 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3453;
        end

       3453 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1151] = 2;
              ip = 3454;
        end

       3454 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[497];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1151];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3455;
              heapClock = 1;
        end

       3455 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3456;
        end

       3456 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1152] = localMem[502];
              ip = 3457;
        end

       3457 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[497];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1152];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 3458;
              heapClock = 1;
        end

       3458 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3459;
        end

       3459 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3527;
        end

       3460 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3461;
        end

       3461 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[498];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3462;
              heapClock = 1;
        end

       3462 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3463;
        end

       3463 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1153] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3464;
              heapClock = 1;
        end

       3464 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3465;
        end

       3465 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[504] = localMem[1153];
              ip = 3466;
        end

       3466 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[504];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[502];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3467;
              heapClock = 1;
        end

       3467 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3468;
        end

       3468 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1154] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3469;
              heapClock = 1;
        end

       3469 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3470;
        end

       3470 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[505] = localMem[1154];
              ip = 3471;
        end

       3471 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[498] = localMem[505];
              ip = 3472;
        end

       3472 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3520;
        end

       3473 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3473");
        end

       3474 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  3474");
        end

       3475 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3475");
        end

       3476 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3476");
        end

       3477 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  3477");
        end

       3478 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3478");
        end

       3479 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3479");
        end

       3480 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3480");
        end

       3481 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3481");
        end

       3482 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3482");
        end

       3483 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3483");
        end

       3484 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  3484");
        end

       3485 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3485");
        end

       3486 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3486");
        end

       3487 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3487");
        end

       3488 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3488");
        end

       3489 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed  3489");
        end

       3490 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  3490");
        end

       3491 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3491");
        end

       3492 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3492");
        end

       3493 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3493");
        end

       3494 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3494");
        end

       3495 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3495");
        end

       3496 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  3496");
        end

       3497 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  3497");
        end

       3498 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3498");
        end

       3499 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3499");
        end

       3500 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3500");
        end

       3501 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3501");
        end

       3502 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3502");
        end

       3503 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3503");
        end

       3504 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3504");
        end

       3505 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  3505");
        end

       3506 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3506");
        end

       3507 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  3507");
        end

       3508 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3508");
        end

       3509 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3509");
        end

       3510 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3510");
        end

       3511 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3511");
        end

       3512 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3512");
        end

       3513 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3513");
        end

       3514 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  3514");
        end

       3515 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3515");
        end

       3516 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  3516");
        end

       3517 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
          // $display("Should not be executed  3517");
        end

       3518 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3518");
        end

       3519 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  3519");
        end

       3520 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3521;
        end

       3521 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[499] = localMem[499] + 1;
              ip = 3522;
        end

       3522 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 3426;
        end

       3523 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3523");
        end

       3524 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  3524");
        end

       3525 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3525");
        end

       3526 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  3526");
        end

       3527 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 3528;
        end

       3528 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[497];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 3529;
              heapClock = 1;
        end

       3529 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3530;
        end

       3530 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1164] = heapOut;                                                     // Data retrieved from heap memory
              ip = 3531;
              heapClock = 1;
        end

       3531 :
        begin                                                                   // resetHeapClock
          //$display("AAAA %4d %4d resetHeapClock", steps, ip);
              heapClock = 0;
              ip = 3532;
        end

       3532 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[511] = localMem[1164];
              ip = 3533;
        end

       3533 :
        begin                                                                   // out
          //$display("AAAA %4d %4d out", steps, ip);
              outMem[outMemPos] = localMem[511];
              outMemPos = outMemPos + 1;
              ip = 3534;
        end
      endcase
      success = outMem[0] == 0 && outMem[1] == 2 && outMem[2] == 4 && outMem[3] == 6 && outMem[4] == 8 && outMem[5] == 10 && outMem[6] == 12 && outMem[7] == 14 && outMem[8] == 16 && outMem[9] == 18 && outMem[10] == 20 && outMem[11] == 22 && outMem[12] == 24 && outMem[13] == 26 && outMem[14] == 28 && outMem[15] == 30 && outMem[16] == 32 && outMem[17] == 34 && outMem[18] == 36 && outMem[19] == 38 && outMem[20] == 40 && outMem[21] == 42 && outMem[22] == 44 && outMem[23] == 46 && outMem[24] == 48 && outMem[25] == 50 && outMem[26] == 52 && outMem[27] == 54 && outMem[28] == 56 && outMem[29] == 58 && outMem[30] == 60 && outMem[31] == 62 && outMem[32] == 64 && outMem[33] == 66 && outMem[34] == 68 && outMem[35] == 70 && outMem[36] == 72 && outMem[37] == 74 && outMem[38] == 76 && outMem[39] == 78 && outMem[40] == 80 && outMem[41] == 82 && outMem[42] == 84 && outMem[43] == 86 && outMem[44] == 88 && outMem[45] == 90 && outMem[46] == 92 && outMem[47] == 94 && outMem[48] == 96 && outMem[49] == 98 && outMem[50] == 100 && outMem[51] == 102 && outMem[52] == 104 && outMem[53] == 106 && outMem[54] == 108 && outMem[55] == 110 && outMem[56] == 112 && outMem[57] == 114 && outMem[58] == 116 && outMem[59] == 118 && outMem[60] == 120 && outMem[61] == 122 && outMem[62] == 124 && outMem[63] == 126 && outMem[64] == 128 && outMem[65] == 130 && outMem[66] == 2;
      steps = steps + 1;
      finished = steps >  51348;
    end
  end

endmodule
