// Check double frees, over allocation
// Check access to unallocated arrays or elements
// Check push overflow, pop underflow
// Next Message 10000280
`define Reset        1  /* Zero all memory sizes                               */
`define Write        2  /* Write an element                                    */
`define Read         3  /* Read an element                                     */
`define Size         4  /* Size of array                                       */
`define Inc          5  /* Increment size of array if possible                 */
`define Dec          6  /* Decrement size of array if possible                 */
`define Index        7  /* Index of element in array                           */
`define Less         8  /* Elements of array less than in                      */
`define Greater      9  /* Elements of array greater than in                   */
`define Up          10  /* Move array up                                       */
`define Down        11  /* Move array down                                     */
`define Long1       12  /* Move long first step                                */
`define Long2       13  /* Move long last  step                                */
`define Push        14  /* Push if possible                                    */
`define Pop         15  /* Pop if possible                                     */
`define Dump        16  /* Dump                                                */
`define Resize      17  /* Resize an array                                     */
`define Alloc       18  /* Allocate a new array before using it                */
`define Free        19  /* Free an array for reuse                             */
`define Add         20  /* Add to an element returning the new value           */
`define AddAfter    21  /* Add to an element returning the previous value      */
`define Subtract    22  /* Subtract to an element returning the new value      */
`define SubAfter    23  /* Subtract to an element returning the previous value */
`define ShiftLeft   24  /* Shift left                                          */
`define ShiftRight  25  /* Shift right                                         */
`define NotLogical  26  /* Not - logical                                       */
`define Not         27  /* Not - bitwise                                       */
`define Or          28  /* Or                                                  */
`define Xor         29  /* Xor                                                 */
`define And         30  /* And                                                 */

module Memory
#(parameter integer ADDRESS_BITS =  8,                                          // Number of bits in an address
  parameter integer INDEX_BITS   =  3,                                          // Bits in in an index
  parameter integer DATA_BITS    = 16)                                          // Width of an element in bits
 (input wire                    clock,                                          // Clock to drive array operations
  input wire[7:0]               action,                                         // Operation to be performed on array
  input wire [ADDRESS_BITS-1:0] array,                                          // The number of the array to work on
  input wire [INDEX_BITS  -1:0] index,                                          // Index within array
  input wire [DATA_BITS   -1:0] in,                                             // Input data
  output reg [DATA_BITS   -1:0] out,                                            // Output data
  output reg [31:0]             error);                                         // Error

  parameter integer ARRAY_LENGTH = 2**INDEX_BITS;                               // Maximum index
  parameter integer ARRAYS       = 2**ADDRESS_BITS;                             // Number of memory elements for both arrays and elements

  reg [DATA_BITS   -1:0] memory     [ARRAYS-1:0][ARRAY_LENGTH-1:0];             // Memory containing arrays in fixed blocks
  reg [DATA_BITS   -1:0] copy                   [ARRAY_LENGTH-1:0];             // Copy of one array
  reg [INDEX_BITS    :0] arraySizes [ARRAYS-1:0];                               // Current size of each array
  reg [ADDRESS_BITS-1:0] freedArrays[ARRAYS-1:0];                               // Currently freed arrays
  reg                    allocations[ARRAYS-1:0];                               // Currently allocated arrays

  integer allocatedArrays;                                                      // Arrays allocated
  integer freedArraysTop;                                                       // Top of the freed arrays stack
  integer result;                                                               // Result of each array operation
  integer size;                                                                 // Size of current array
  integer moveLongStartArray;                                                   // Source array of move long
  integer moveLongStartIndex;                                                   // Source index of move long
  integer i, a, b;                                                              // Index

  task checkWriteable(input integer err);                                       // Check a memory is writable
    begin
       error = 0;
       if (array >= allocatedArrays) begin
         //$display("Array has not been allocated, array %d", array);
         error = err;
       end
       if (!allocations[array]) begin
         //$display("Array has been freed, array %d", array);
         error = err + 1;
       end
    end
  endtask

  task checkReadable(input integer err);                                        // Check a memory locationis readable
    begin
       checkWriteable(err);
       if (index >= arraySizes[array]) begin
         //$display("Access outside array bounds, array %d, size: %d, access: %d", array, arraySizes[array], index);
         error = err + 2;
       end
    end
  endtask

  task dump;                                                                    // Dump some memory
    begin
      //$display("    %2d %2d %2d", arraySizes[0], arraySizes[1], arraySizes[2]);
      for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
        //$display("%2d  %2d %2d %2d", i, memory[0][i], memory[1][i], memory[2][i]);
      end
    end
  endtask

  always @(clock) begin                                                             // Each transition
    case(action)                                                                // Decode request
      `Reset: begin                                                             // Reset
        freedArraysTop = 0;                                                     // Free all arrays
        allocatedArrays = 0;
      end

      `Write: begin                                                             // Write
        checkWriteable(10000010);
        if (!error) begin
          memory[array][index] = in;
          if (index >= arraySizes[array] && index < ARRAY_LENGTH) begin
            arraySizes[array] = index + 1;
          end
          out = in;
        end
      end

      `Read: begin                                                              // Read
        checkReadable(10000020);
        if (!error) begin
          out = memory[array][index];
        end
      end

      `Size: begin                                                              // Size
        checkWriteable(10000030);
        if (!error) begin
          out = arraySizes[array];
        end
      end

      `Dec: begin                                                               // Decrement
        checkWriteable(10000040);
        if (!error) begin
          if (arraySizes[array] > 0) arraySizes[array] = arraySizes[array] - 1;
          else begin
            //$display("Attempt to decrement empty array, array %d", array); error = 10000044;
          end
        end
      end

      `Inc: begin                                                               // Increment
        checkWriteable(10000050);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;
          else begin
            //$display("Attempt to decrement full array, array %d", array);  error = 10000054;
          end
        end
      end

      `Index: begin                                                             // Index
        checkWriteable(10000060);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] == in) result = i + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Less: begin                                                              // Count less
        checkWriteable(10000070);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] < in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Greater: begin                                                           // Count greater
        checkWriteable(10000080);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] > in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Down: begin                                                              // Down
        checkWriteable(10000270);
        if (!error) begin
          size   = arraySizes[array];
          if (size > 0) begin
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i]; // Copy source array
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                       // Move original array up
              if (i > index && i <= size) begin
                memory[array][i-1] = copy[i];
              end
            end
            out = copy[index];                                                  // Return replaced value
            arraySizes[array] = arraySizes[array] - 1;                          // Decrease array size
          end
          else error = 100000274;                                               // Orignal array was emoty so we cannot shift it down
        end
      end

      `Up: begin                                                                // Up
        checkWriteable(10000090);
        if (!error) begin
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i];   // Copy source array
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Move original array up
            if (i > index && i <= size) begin
              memory[array][i] = copy[i-1];
            end
          end
          memory[array][index] = in;                                            // Insert new value
          if (size < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;   // Increase array size
        end
      end

      `Long1: begin                                                             // Move long start
        checkReadable(10000100);
        if (!error) begin
          moveLongStartArray = array;                                           // Record source
          moveLongStartIndex = index;
        end
      end

      `Long2: begin                                                             // Move long finish
        checkWriteable(10000110);
        if (!error) begin
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Copy from source to target
            if (i < in && index + i < ARRAY_LENGTH && moveLongStartIndex+i < ARRAY_LENGTH) begin
              memory[array][index+i] = memory[moveLongStartArray][moveLongStartIndex+i];
              if (index+i >= arraySizes[array]) arraySizes[array] = index+i+1;
            end
          end
        end
      end

      `Push: begin                                                              // Push
        checkWriteable(10000120);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) begin
            memory[array][arraySizes[array]] = in;
            arraySizes[array] = arraySizes[array] + 1;
          end
          else begin
            //$display("Attempt to push to full array, array %d, value %d", array, in);  error = 10000124;
          end
        end
      end

      `Pop: begin                                                               // Pop
        checkWriteable(10000130);
        if (!error) begin
          if (arraySizes[array] > 0) begin
            arraySizes[array] = arraySizes[array] - 1;
            out = memory[array][arraySizes[array]];
          end
          else begin
            //$display("Attempt to pop empty array, array %d", array); error = 10000134;
          end
        end
      end

      `Dump: begin                                                              // Dump
        dump();
      end

      `Resize: begin                                                            // Resize
        checkWriteable(10000140);
        if (!error) begin
          if (in <= ARRAY_LENGTH) arraySizes[array] = in;
          else begin
            //$display("Attempt to make an array too large, array %d, max %d, size %d", array, ARRAY_LENGTH, in); error = 10000144;
          end
        end
      end

      `Alloc: begin                                                             // Allocate an array
        if (freedArraysTop > 0) begin                                           // Reuse a freed array
          freedArraysTop = freedArraysTop - 1;
          result = freedArrays[freedArraysTop];
        end
        else if (allocatedArrays < ARRAYS-1) begin                              // Allocate a new array - assumes enough memory
          result          = allocatedArrays;
          allocatedArrays = allocatedArrays + 1;
        end
        else begin
          //$display("Out of memory, cannot allocate a new array"); error = 10000270;
        end
        allocations[result] = 1;                                                // Allocated
        arraySizes[result] = 0;                                                 // Empty array
        out = result;
      end

      `Free: begin                                                              // Free an array
        checkWriteable(10000150);
        if (!error) begin
          freedArrays[freedArraysTop] = array;                                  // Relies on the user not re freeing a freed array - we should probably hve another array to prevent this
          allocations[freedArraysTop] = 0;                                      // No longer allocated
          freedArraysTop = freedArraysTop + 1;
        end
      end

      `Add: begin                                                               // Add to an element
        checkReadable(10000160);
        if (!error) begin
          memory[array][index] = memory[array][index] + in;
          out = memory[array][index];
        end
      end

      `AddAfter: begin                                                          // Add to an element after putting the content of the element on out
        checkReadable(10000170);
        if (!error) begin
        out = memory[array][index];
        memory[array][index] = memory[array][index] + in;
        end
      end

      `Subtract: begin                                                          // Subtract from an element
        checkReadable(10000180);
        if (!error) begin
          memory[array][index] = memory[array][index] - in;
          out = memory[array][index];
        end
      end

      `SubAfter: begin                                                          // Subtract from an element after putting the content of the element on out
        checkReadable(10000190);
        if (!error) begin
          out = memory[array][index];
          memory[array][index] = memory[array][index] - in;
        end
      end

      `ShiftLeft: begin                                                         // Shift left
        checkReadable(10000200);
        if (!error) begin
          memory[array][index] = memory[array][index] << in;
          out = memory[array][index];
        end
      end

      `ShiftRight: begin                                                        // Shift right
        checkReadable(10000210);
        if (!error) begin
          memory[array][index] = memory[array][index] >> in;
          out = memory[array][index];
        end
      end

      `NotLogical: begin                                                        // Not logical
        checkReadable(10000220);
        if (!error) begin
          memory[array][index] = !memory[array][index];
          out = memory[array][index];
        end
      end

      `Not: begin                                                               // Not
        checkReadable(10000230);
        if (!error) begin
          memory[array][index] = ~memory[array][index];
          out = memory[array][index];
        end
      end

      `Or: begin                                                                // Or
        checkReadable(10000240);
        if (!error) begin
          memory[array][index] = memory[array][index] | in;
          out = memory[array][index];
        end
      end

      `Xor: begin                                                               // Xor
        checkReadable(10000250);
        if (!error) begin
          memory[array][index] = memory[array][index] ^ in;
          out = memory[array][index];
        end
      end

      `And: begin                                                               // And
        checkReadable(10000260);
        if (!error) begin
          memory[array][index] = memory[array][index] & in;
          out = memory[array][index];
        end
      end
    endcase
  end
endmodule
//-----------------------------------------------------------------------------
// Fpga test
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga                                                                     // Run test programs
 (input  wire clock,                                                            // Driving clock
  input  wire reset,                                                            // Restart program
  output reg  finished,                                                         // Goes high when the program has finished
  output reg  success);                                                         // Goes high on finish if all the tests passed

  reg                heapClock;                                                 // Clock to drive array operations
  reg [7:0]          heapAction;                                                // Operation to be performed on array
  reg [       3-1:0] heapArray;                                         // The number of the array to work on
  reg [       3-1:0] heapIndex;                                         // Index within array
  reg [      12-1:0] heapIn;                                            // Input data
  reg [      12-1:0] heapOut;                                           // Output data
  reg [31        :0] heapError;                                                 // Error on heap operation if not zero

  Memory                                                                        // Memory module
   #(       3,        3,       12)                          // Address bits, index bits, data bits
    heap(                                                                       // Create heap memory
    .clock  (heapClock),
    .action (heapAction),
    .array  (heapArray),
    .index  (heapIndex),
    .in     (heapIn),
    .out    (heapOut),
    .error  (heapError)
  );
  reg [      12-1:0] localMem[     500-1:0];                       // Local memory
  reg [      12-1:0]   outMem[       1  -1:0];                       // Out channel
  reg [      12-1:0]    inMem[       1   -1:0];                       // In channel

  integer inMemPos;                                                             // Current position in input channel
  integer outMemPos;                                                            // Position in output channel

  integer ip;                                                                   // Instruction pointer
  integer steps;                                                                // Number of steps executed so far
  integer i, j, k;                                                              // A useful counter

  always @(posedge clock, negedge clock) begin                                  // Each instruction
    if (reset) begin
      ip             = 0;
      steps          = 0;
      inMemPos       = 0;
      outMemPos      = 0;
      finished       = 0;
      success        = 0;

    end
    else begin
      steps = steps + 1;
      case(ip)

          0 :
        begin                                                                   // start
          //$display("AAAA %4d %4d start", steps, ip);
              heapClock = 0;                                                    // Ready for next operation
              ip = 1;
        end

          1 :
        begin                                                                   // start2
          //$display("AAAA %4d %4d start2", steps, ip);
              heapAction = `Reset;                                          // Ready for next operation
              ip = 2;
              heapClock = ~ heapClock;
        end

          2 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3;
              heapClock = ~ heapClock;
        end

          3 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[0] = heapOut;
              ip = 4;
        end

          4 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[476] = 3;
              ip = 5;
        end

          5 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[476];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 6;
              heapClock = ~ heapClock;
        end

          6 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[477] = 0;
              ip = 7;
        end

          7 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[477];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 8;
              heapClock = ~ heapClock;
        end

          8 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[478] = 0;
              ip = 9;
        end

          9 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[478];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 10;
              heapClock = ~ heapClock;
        end

         10 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[479] = 0;
              ip = 11;
        end

         11 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[479];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 12;
              heapClock = ~ heapClock;
        end

         12 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 13;
              heapClock = ~ heapClock;
        end

         13 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[1] = heapOut;
              ip = 14;
        end

         14 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 15;
        end

         15 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 16;
              heapClock = ~ heapClock;
        end

         16 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[480] = heapOut;                                                     // Data retrieved from heap memory
              ip = 17;
              heapClock = ~ heapClock;
        end

         17 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[2] = localMem[480];
              ip = 18;
        end

         18 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[2] != 0 ? 70 : 19;
        end

         19 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 20;
              heapClock = ~ heapClock;
        end

         20 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[3] = heapOut;
              ip = 21;
        end

         21 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = 1;
              ip = 22;
        end

         22 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[481];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 23;
              heapClock = ~ heapClock;
        end

         23 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[482] = 0;
              ip = 24;
        end

         24 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[482];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 25;
              heapClock = ~ heapClock;
        end

         25 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 26;
              heapClock = ~ heapClock;
        end

         26 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[4] = heapOut;
              ip = 27;
        end

         27 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[483] = localMem[4];
              ip = 28;
        end

         28 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[483];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 29;
              heapClock = ~ heapClock;
        end

         29 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 30;
              heapClock = ~ heapClock;
        end

         30 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[5] = heapOut;
              ip = 31;
        end

         31 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[484] = localMem[5];
              ip = 32;
        end

         32 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[484];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 33;
              heapClock = ~ heapClock;
        end

         33 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[485] = 0;
              ip = 34;
        end

         34 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[485];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 35;
              heapClock = ~ heapClock;
        end

         35 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[486] = localMem[0];
              ip = 36;
        end

         36 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[486];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 37;
              heapClock = ~ heapClock;
        end

         37 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 38;
              heapClock = ~ heapClock;
        end

         38 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[487] = heapOut;                                                     // Data retrieved from heap memory
              ip = 39;
              heapClock = ~ heapClock;
        end

         39 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[488] = localMem[487] + 1;
              ip = 40;
        end

         40 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[488];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 41;
              heapClock = ~ heapClock;
        end

         41 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 42;
              heapClock = ~ heapClock;
        end

         42 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[489] = heapOut;                                                     // Data retrieved from heap memory
              ip = 43;
              heapClock = ~ heapClock;
        end

         43 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[490] = localMem[489];
              ip = 44;
        end

         44 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[3];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[490];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 45;
              heapClock = ~ heapClock;
        end

         45 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 46;
              heapClock = ~ heapClock;
        end

         46 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[491] = heapOut;                                                     // Data retrieved from heap memory
              ip = 47;
              heapClock = ~ heapClock;
        end

         47 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[6] = localMem[491];
              ip = 48;
        end

         48 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[492] = 1;
              ip = 49;
        end

         49 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[6];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[492];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 50;
              heapClock = ~ heapClock;
        end

         50 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 51;
              heapClock = ~ heapClock;
        end

         51 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[493] = heapOut;                                                     // Data retrieved from heap memory
              ip = 52;
              heapClock = ~ heapClock;
        end

         52 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[7] = localMem[493];
              ip = 53;
        end

         53 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[494] = 11;
              ip = 54;
        end

         54 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[494];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 55;
              heapClock = ~ heapClock;
        end

         55 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 56;
              heapClock = ~ heapClock;
        end

         56 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[495] = heapOut;                                                     // Data retrieved from heap memory
              ip = 57;
              heapClock = ~ heapClock;
        end

         57 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[496] = localMem[495] + 1;
              ip = 58;
        end

         58 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[496];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 59;
              heapClock = ~ heapClock;
        end

         59 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[497] = localMem[3];
              ip = 60;
        end

         60 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[497];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 61;
              heapClock = ~ heapClock;
        end

         61 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 62;
              heapClock = ~ heapClock;
        end

         62 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[498] = heapOut;                                                     // Data retrieved from heap memory
              ip = 63;
              heapClock = ~ heapClock;
        end

         63 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[8] = localMem[498];
              ip = 64;
        end

         64 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[8];
              ip = 65;
              heapClock = ~ heapClock;
        end

         65 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[3];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 66;
              heapClock = ~ heapClock;
        end

         66 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[499] = heapOut;                                                     // Data retrieved from heap memory
              ip = 67;
              heapClock = ~ heapClock;
        end

         67 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[9] = localMem[499];
              ip = 68;
        end

         68 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[9];
              ip = 69;
              heapClock = ~ heapClock;
        end

         69 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2179;
        end

         70 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed    70");
        end

         71 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed    71");
        end

         72 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed    72");
        end

         73 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed    73");
        end

         74 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed    74");
        end

         75 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed    75");
        end

         76 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed    76");
        end

         77 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed    77");
        end

         78 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed    78");
        end

         79 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed    79");
        end

         80 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed    80");
        end

         81 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed    81");
        end

         82 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed    82");
        end

         83 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed    83");
        end

         84 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed    84");
        end

         85 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed    85");
        end

         86 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed    86");
        end

         87 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed    87");
        end

         88 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed    88");
        end

         89 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed    89");
        end

         90 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed    90");
        end

         91 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed    91");
        end

         92 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed    92");
        end

         93 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed    93");
        end

         94 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed    94");
        end

         95 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed    95");
        end

         96 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed    96");
        end

         97 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed    97");
        end

         98 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed    98");
        end

         99 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed    99");
        end

        100 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   100");
        end

        101 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   101");
        end

        102 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   102");
        end

        103 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   103");
        end

        104 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   104");
        end

        105 :
        begin                                                                   // arrayCountGreater
          //$display("AAAA %4d %4d arrayCountGreater", steps, ip);
          // $display("Should not be executed   105");
        end

        106 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   106");
        end

        107 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   107");
        end

        108 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   108");
        end

        109 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   109");
        end

        110 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   110");
        end

        111 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   111");
        end

        112 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   112");
        end

        113 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   113");
        end

        114 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   114");
        end

        115 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   115");
        end

        116 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   116");
        end

        117 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   117");
        end

        118 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   118");
        end

        119 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   119");
        end

        120 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   120");
        end

        121 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   121");
        end

        122 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   122");
        end

        123 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   123");
        end

        124 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   124");
        end

        125 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   125");
        end

        126 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed   126");
        end

        127 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   127");
        end

        128 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   128");
        end

        129 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   129");
        end

        130 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   130");
        end

        131 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   131");
        end

        132 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   132");
        end

        133 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   133");
        end

        134 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   134");
        end

        135 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   135");
        end

        136 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   136");
        end

        137 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   137");
        end

        138 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   138");
        end

        139 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   139");
        end

        140 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   140");
        end

        141 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   141");
        end

        142 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   142");
        end

        143 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   143");
        end

        144 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   144");
        end

        145 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   145");
        end

        146 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   146");
        end

        147 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   147");
        end

        148 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   148");
        end

        149 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   149");
        end

        150 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   150");
        end

        151 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   151");
        end

        152 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   152");
        end

        153 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   153");
        end

        154 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   154");
        end

        155 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   155");
        end

        156 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   156");
        end

        157 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   157");
        end

        158 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   158");
        end

        159 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   159");
        end

        160 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   160");
        end

        161 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
          // $display("Should not be executed   161");
        end

        162 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   162");
        end

        163 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
          // $display("Should not be executed   163");
        end

        164 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   164");
        end

        165 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   165");
        end

        166 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   166");
        end

        167 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   167");
        end

        168 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed   168");
        end

        169 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   169");
        end

        170 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   170");
        end

        171 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   171");
        end

        172 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   172");
        end

        173 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   173");
        end

        174 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   174");
        end

        175 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   175");
        end

        176 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   176");
        end

        177 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   177");
        end

        178 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   178");
        end

        179 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   179");
        end

        180 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   180");
        end

        181 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   181");
        end

        182 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   182");
        end

        183 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   183");
        end

        184 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   184");
        end

        185 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   185");
        end

        186 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   186");
        end

        187 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   187");
        end

        188 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   188");
        end

        189 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   189");
        end

        190 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   190");
        end

        191 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   191");
        end

        192 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   192");
        end

        193 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   193");
        end

        194 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   194");
        end

        195 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   195");
        end

        196 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   196");
        end

        197 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   197");
        end

        198 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   198");
        end

        199 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   199");
        end

        200 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   200");
        end

        201 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   201");
        end

        202 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   202");
        end

        203 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   203");
        end

        204 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   204");
        end

        205 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   205");
        end

        206 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   206");
        end

        207 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   207");
        end

        208 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   208");
        end

        209 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   209");
        end

        210 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   210");
        end

        211 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   211");
        end

        212 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   212");
        end

        213 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   213");
        end

        214 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   214");
        end

        215 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   215");
        end

        216 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   216");
        end

        217 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   217");
        end

        218 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   218");
        end

        219 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   219");
        end

        220 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   220");
        end

        221 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   221");
        end

        222 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   222");
        end

        223 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   223");
        end

        224 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   224");
        end

        225 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   225");
        end

        226 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   226");
        end

        227 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   227");
        end

        228 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   228");
        end

        229 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   229");
        end

        230 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   230");
        end

        231 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   231");
        end

        232 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   232");
        end

        233 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   233");
        end

        234 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   234");
        end

        235 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   235");
        end

        236 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   236");
        end

        237 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   237");
        end

        238 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   238");
        end

        239 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   239");
        end

        240 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   240");
        end

        241 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   241");
        end

        242 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   242");
        end

        243 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   243");
        end

        244 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   244");
        end

        245 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   245");
        end

        246 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   246");
        end

        247 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   247");
        end

        248 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   248");
        end

        249 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   249");
        end

        250 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   250");
        end

        251 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   251");
        end

        252 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   252");
        end

        253 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   253");
        end

        254 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   254");
        end

        255 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   255");
        end

        256 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   256");
        end

        257 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   257");
        end

        258 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   258");
        end

        259 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   259");
        end

        260 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   260");
        end

        261 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   261");
        end

        262 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   262");
        end

        263 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   263");
        end

        264 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   264");
        end

        265 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   265");
        end

        266 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   266");
        end

        267 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   267");
        end

        268 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   268");
        end

        269 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   269");
        end

        270 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   270");
        end

        271 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   271");
        end

        272 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   272");
        end

        273 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   273");
        end

        274 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   274");
        end

        275 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   275");
        end

        276 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   276");
        end

        277 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   277");
        end

        278 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   278");
        end

        279 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   279");
        end

        280 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   280");
        end

        281 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   281");
        end

        282 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   282");
        end

        283 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   283");
        end

        284 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   284");
        end

        285 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   285");
        end

        286 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   286");
        end

        287 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   287");
        end

        288 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   288");
        end

        289 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   289");
        end

        290 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   290");
        end

        291 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   291");
        end

        292 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   292");
        end

        293 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   293");
        end

        294 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   294");
        end

        295 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   295");
        end

        296 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   296");
        end

        297 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   297");
        end

        298 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   298");
        end

        299 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   299");
        end

        300 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   300");
        end

        301 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   301");
        end

        302 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   302");
        end

        303 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   303");
        end

        304 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   304");
        end

        305 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   305");
        end

        306 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   306");
        end

        307 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   307");
        end

        308 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   308");
        end

        309 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   309");
        end

        310 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   310");
        end

        311 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   311");
        end

        312 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   312");
        end

        313 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   313");
        end

        314 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   314");
        end

        315 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   315");
        end

        316 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   316");
        end

        317 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   317");
        end

        318 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   318");
        end

        319 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   319");
        end

        320 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   320");
        end

        321 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   321");
        end

        322 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   322");
        end

        323 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   323");
        end

        324 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   324");
        end

        325 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   325");
        end

        326 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   326");
        end

        327 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   327");
        end

        328 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   328");
        end

        329 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   329");
        end

        330 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   330");
        end

        331 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   331");
        end

        332 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   332");
        end

        333 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   333");
        end

        334 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   334");
        end

        335 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   335");
        end

        336 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   336");
        end

        337 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   337");
        end

        338 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   338");
        end

        339 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   339");
        end

        340 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   340");
        end

        341 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   341");
        end

        342 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   342");
        end

        343 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   343");
        end

        344 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   344");
        end

        345 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   345");
        end

        346 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   346");
        end

        347 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   347");
        end

        348 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   348");
        end

        349 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   349");
        end

        350 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   350");
        end

        351 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   351");
        end

        352 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   352");
        end

        353 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   353");
        end

        354 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   354");
        end

        355 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   355");
        end

        356 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   356");
        end

        357 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   357");
        end

        358 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   358");
        end

        359 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   359");
        end

        360 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   360");
        end

        361 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   361");
        end

        362 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   362");
        end

        363 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   363");
        end

        364 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   364");
        end

        365 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   365");
        end

        366 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   366");
        end

        367 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   367");
        end

        368 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   368");
        end

        369 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   369");
        end

        370 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   370");
        end

        371 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   371");
        end

        372 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   372");
        end

        373 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   373");
        end

        374 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   374");
        end

        375 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   375");
        end

        376 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   376");
        end

        377 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   377");
        end

        378 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   378");
        end

        379 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   379");
        end

        380 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   380");
        end

        381 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   381");
        end

        382 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   382");
        end

        383 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   383");
        end

        384 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   384");
        end

        385 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   385");
        end

        386 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   386");
        end

        387 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   387");
        end

        388 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   388");
        end

        389 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   389");
        end

        390 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   390");
        end

        391 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   391");
        end

        392 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   392");
        end

        393 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   393");
        end

        394 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   394");
        end

        395 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   395");
        end

        396 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   396");
        end

        397 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   397");
        end

        398 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   398");
        end

        399 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   399");
        end

        400 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   400");
        end

        401 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   401");
        end

        402 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   402");
        end

        403 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   403");
        end

        404 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   404");
        end

        405 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   405");
        end

        406 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   406");
        end

        407 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   407");
        end

        408 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   408");
        end

        409 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   409");
        end

        410 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   410");
        end

        411 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   411");
        end

        412 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   412");
        end

        413 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   413");
        end

        414 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   414");
        end

        415 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   415");
        end

        416 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   416");
        end

        417 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   417");
        end

        418 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   418");
        end

        419 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   419");
        end

        420 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   420");
        end

        421 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   421");
        end

        422 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   422");
        end

        423 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   423");
        end

        424 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   424");
        end

        425 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   425");
        end

        426 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   426");
        end

        427 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   427");
        end

        428 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   428");
        end

        429 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   429");
        end

        430 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   430");
        end

        431 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   431");
        end

        432 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   432");
        end

        433 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   433");
        end

        434 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   434");
        end

        435 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   435");
        end

        436 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   436");
        end

        437 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   437");
        end

        438 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   438");
        end

        439 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   439");
        end

        440 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   440");
        end

        441 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   441");
        end

        442 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   442");
        end

        443 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   443");
        end

        444 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   444");
        end

        445 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   445");
        end

        446 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   446");
        end

        447 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   447");
        end

        448 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   448");
        end

        449 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   449");
        end

        450 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   450");
        end

        451 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   451");
        end

        452 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   452");
        end

        453 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   453");
        end

        454 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   454");
        end

        455 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   455");
        end

        456 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   456");
        end

        457 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   457");
        end

        458 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   458");
        end

        459 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   459");
        end

        460 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   460");
        end

        461 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   461");
        end

        462 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   462");
        end

        463 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   463");
        end

        464 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   464");
        end

        465 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   465");
        end

        466 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   466");
        end

        467 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   467");
        end

        468 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   468");
        end

        469 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   469");
        end

        470 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   470");
        end

        471 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   471");
        end

        472 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   472");
        end

        473 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   473");
        end

        474 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   474");
        end

        475 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   475");
        end

        476 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   476");
        end

        477 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   477");
        end

        478 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   478");
        end

        479 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   479");
        end

        480 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   480");
        end

        481 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   481");
        end

        482 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   482");
        end

        483 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   483");
        end

        484 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   484");
        end

        485 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   485");
        end

        486 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   486");
        end

        487 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   487");
        end

        488 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   488");
        end

        489 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   489");
        end

        490 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   490");
        end

        491 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   491");
        end

        492 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   492");
        end

        493 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   493");
        end

        494 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   494");
        end

        495 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   495");
        end

        496 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   496");
        end

        497 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   497");
        end

        498 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   498");
        end

        499 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   499");
        end

        500 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   500");
        end

        501 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   501");
        end

        502 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   502");
        end

        503 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   503");
        end

        504 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   504");
        end

        505 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   505");
        end

        506 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   506");
        end

        507 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   507");
        end

        508 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   508");
        end

        509 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   509");
        end

        510 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   510");
        end

        511 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   511");
        end

        512 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   512");
        end

        513 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   513");
        end

        514 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   514");
        end

        515 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   515");
        end

        516 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   516");
        end

        517 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   517");
        end

        518 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   518");
        end

        519 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   519");
        end

        520 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   520");
        end

        521 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   521");
        end

        522 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   522");
        end

        523 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   523");
        end

        524 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   524");
        end

        525 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   525");
        end

        526 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   526");
        end

        527 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   527");
        end

        528 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   528");
        end

        529 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   529");
        end

        530 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   530");
        end

        531 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   531");
        end

        532 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   532");
        end

        533 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   533");
        end

        534 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   534");
        end

        535 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   535");
        end

        536 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   536");
        end

        537 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   537");
        end

        538 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   538");
        end

        539 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   539");
        end

        540 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   540");
        end

        541 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   541");
        end

        542 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   542");
        end

        543 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   543");
        end

        544 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   544");
        end

        545 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   545");
        end

        546 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   546");
        end

        547 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   547");
        end

        548 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   548");
        end

        549 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   549");
        end

        550 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   550");
        end

        551 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   551");
        end

        552 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   552");
        end

        553 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   553");
        end

        554 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   554");
        end

        555 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   555");
        end

        556 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   556");
        end

        557 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   557");
        end

        558 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   558");
        end

        559 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   559");
        end

        560 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   560");
        end

        561 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   561");
        end

        562 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   562");
        end

        563 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   563");
        end

        564 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   564");
        end

        565 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   565");
        end

        566 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   566");
        end

        567 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   567");
        end

        568 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   568");
        end

        569 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   569");
        end

        570 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   570");
        end

        571 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   571");
        end

        572 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   572");
        end

        573 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   573");
        end

        574 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   574");
        end

        575 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   575");
        end

        576 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   576");
        end

        577 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   577");
        end

        578 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   578");
        end

        579 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   579");
        end

        580 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   580");
        end

        581 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   581");
        end

        582 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   582");
        end

        583 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   583");
        end

        584 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   584");
        end

        585 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   585");
        end

        586 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   586");
        end

        587 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   587");
        end

        588 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   588");
        end

        589 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   589");
        end

        590 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   590");
        end

        591 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   591");
        end

        592 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   592");
        end

        593 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   593");
        end

        594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   594");
        end

        595 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   595");
        end

        596 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   596");
        end

        597 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   597");
        end

        598 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   598");
        end

        599 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   599");
        end

        600 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   600");
        end

        601 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   601");
        end

        602 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   602");
        end

        603 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   603");
        end

        604 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   604");
        end

        605 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   605");
        end

        606 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   606");
        end

        607 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   607");
        end

        608 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   608");
        end

        609 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   609");
        end

        610 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   610");
        end

        611 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   611");
        end

        612 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   612");
        end

        613 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   613");
        end

        614 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   614");
        end

        615 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   615");
        end

        616 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   616");
        end

        617 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   617");
        end

        618 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   618");
        end

        619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   619");
        end

        620 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   620");
        end

        621 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   621");
        end

        622 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   622");
        end

        623 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   623");
        end

        624 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   624");
        end

        625 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   625");
        end

        626 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   626");
        end

        627 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   627");
        end

        628 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   628");
        end

        629 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   629");
        end

        630 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   630");
        end

        631 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   631");
        end

        632 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   632");
        end

        633 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   633");
        end

        634 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   634");
        end

        635 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   635");
        end

        636 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   636");
        end

        637 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   637");
        end

        638 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   638");
        end

        639 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
          // $display("Should not be executed   639");
        end

        640 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   640");
        end

        641 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   641");
        end

        642 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   642");
        end

        643 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed   643");
        end

        644 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   644");
        end

        645 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   645");
        end

        646 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   646");
        end

        647 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   647");
        end

        648 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   648");
        end

        649 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   649");
        end

        650 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   650");
        end

        651 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   651");
        end

        652 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   652");
        end

        653 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   653");
        end

        654 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   654");
        end

        655 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   655");
        end

        656 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   656");
        end

        657 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   657");
        end

        658 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   658");
        end

        659 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   659");
        end

        660 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   660");
        end

        661 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   661");
        end

        662 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   662");
        end

        663 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   663");
        end

        664 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   664");
        end

        665 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   665");
        end

        666 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   666");
        end

        667 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   667");
        end

        668 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
          // $display("Should not be executed   668");
        end

        669 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   669");
        end

        670 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
          // $display("Should not be executed   670");
        end

        671 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   671");
        end

        672 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   672");
        end

        673 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   673");
        end

        674 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   674");
        end

        675 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed   675");
        end

        676 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   676");
        end

        677 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   677");
        end

        678 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   678");
        end

        679 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   679");
        end

        680 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   680");
        end

        681 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   681");
        end

        682 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   682");
        end

        683 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   683");
        end

        684 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   684");
        end

        685 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   685");
        end

        686 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   686");
        end

        687 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   687");
        end

        688 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   688");
        end

        689 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   689");
        end

        690 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   690");
        end

        691 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   691");
        end

        692 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   692");
        end

        693 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   693");
        end

        694 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   694");
        end

        695 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   695");
        end

        696 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   696");
        end

        697 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   697");
        end

        698 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   698");
        end

        699 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   699");
        end

        700 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   700");
        end

        701 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   701");
        end

        702 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   702");
        end

        703 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   703");
        end

        704 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   704");
        end

        705 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   705");
        end

        706 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   706");
        end

        707 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   707");
        end

        708 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   708");
        end

        709 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   709");
        end

        710 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   710");
        end

        711 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   711");
        end

        712 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   712");
        end

        713 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   713");
        end

        714 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   714");
        end

        715 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   715");
        end

        716 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   716");
        end

        717 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   717");
        end

        718 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   718");
        end

        719 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   719");
        end

        720 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   720");
        end

        721 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   721");
        end

        722 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   722");
        end

        723 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   723");
        end

        724 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   724");
        end

        725 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   725");
        end

        726 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   726");
        end

        727 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   727");
        end

        728 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   728");
        end

        729 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   729");
        end

        730 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   730");
        end

        731 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   731");
        end

        732 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   732");
        end

        733 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   733");
        end

        734 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   734");
        end

        735 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   735");
        end

        736 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   736");
        end

        737 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   737");
        end

        738 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   738");
        end

        739 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   739");
        end

        740 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   740");
        end

        741 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   741");
        end

        742 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   742");
        end

        743 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   743");
        end

        744 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   744");
        end

        745 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   745");
        end

        746 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   746");
        end

        747 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   747");
        end

        748 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   748");
        end

        749 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   749");
        end

        750 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   750");
        end

        751 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   751");
        end

        752 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   752");
        end

        753 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   753");
        end

        754 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   754");
        end

        755 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   755");
        end

        756 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   756");
        end

        757 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   757");
        end

        758 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   758");
        end

        759 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   759");
        end

        760 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   760");
        end

        761 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   761");
        end

        762 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   762");
        end

        763 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   763");
        end

        764 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   764");
        end

        765 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   765");
        end

        766 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   766");
        end

        767 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   767");
        end

        768 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   768");
        end

        769 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   769");
        end

        770 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   770");
        end

        771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   771");
        end

        772 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   772");
        end

        773 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   773");
        end

        774 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   774");
        end

        775 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   775");
        end

        776 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   776");
        end

        777 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   777");
        end

        778 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   778");
        end

        779 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   779");
        end

        780 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   780");
        end

        781 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   781");
        end

        782 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   782");
        end

        783 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   783");
        end

        784 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   784");
        end

        785 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   785");
        end

        786 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   786");
        end

        787 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   787");
        end

        788 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   788");
        end

        789 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   789");
        end

        790 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   790");
        end

        791 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   791");
        end

        792 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   792");
        end

        793 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   793");
        end

        794 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   794");
        end

        795 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   795");
        end

        796 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   796");
        end

        797 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   797");
        end

        798 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   798");
        end

        799 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   799");
        end

        800 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   800");
        end

        801 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   801");
        end

        802 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   802");
        end

        803 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   803");
        end

        804 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   804");
        end

        805 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   805");
        end

        806 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   806");
        end

        807 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   807");
        end

        808 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   808");
        end

        809 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   809");
        end

        810 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   810");
        end

        811 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   811");
        end

        812 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   812");
        end

        813 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   813");
        end

        814 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   814");
        end

        815 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   815");
        end

        816 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   816");
        end

        817 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   817");
        end

        818 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   818");
        end

        819 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   819");
        end

        820 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   820");
        end

        821 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   821");
        end

        822 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   822");
        end

        823 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   823");
        end

        824 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   824");
        end

        825 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   825");
        end

        826 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   826");
        end

        827 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   827");
        end

        828 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   828");
        end

        829 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   829");
        end

        830 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   830");
        end

        831 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   831");
        end

        832 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   832");
        end

        833 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   833");
        end

        834 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   834");
        end

        835 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   835");
        end

        836 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   836");
        end

        837 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   837");
        end

        838 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   838");
        end

        839 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   839");
        end

        840 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   840");
        end

        841 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   841");
        end

        842 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   842");
        end

        843 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   843");
        end

        844 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   844");
        end

        845 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   845");
        end

        846 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   846");
        end

        847 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   847");
        end

        848 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   848");
        end

        849 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   849");
        end

        850 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   850");
        end

        851 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   851");
        end

        852 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   852");
        end

        853 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   853");
        end

        854 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   854");
        end

        855 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   855");
        end

        856 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   856");
        end

        857 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   857");
        end

        858 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   858");
        end

        859 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   859");
        end

        860 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   860");
        end

        861 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   861");
        end

        862 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   862");
        end

        863 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   863");
        end

        864 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   864");
        end

        865 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   865");
        end

        866 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   866");
        end

        867 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   867");
        end

        868 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   868");
        end

        869 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   869");
        end

        870 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   870");
        end

        871 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   871");
        end

        872 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   872");
        end

        873 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   873");
        end

        874 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   874");
        end

        875 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   875");
        end

        876 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   876");
        end

        877 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   877");
        end

        878 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   878");
        end

        879 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   879");
        end

        880 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   880");
        end

        881 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   881");
        end

        882 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   882");
        end

        883 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   883");
        end

        884 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   884");
        end

        885 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   885");
        end

        886 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   886");
        end

        887 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   887");
        end

        888 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   888");
        end

        889 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   889");
        end

        890 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   890");
        end

        891 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   891");
        end

        892 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   892");
        end

        893 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   893");
        end

        894 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   894");
        end

        895 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   895");
        end

        896 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   896");
        end

        897 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   897");
        end

        898 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   898");
        end

        899 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   899");
        end

        900 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   900");
        end

        901 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   901");
        end

        902 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   902");
        end

        903 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   903");
        end

        904 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   904");
        end

        905 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   905");
        end

        906 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   906");
        end

        907 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   907");
        end

        908 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   908");
        end

        909 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   909");
        end

        910 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   910");
        end

        911 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   911");
        end

        912 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   912");
        end

        913 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   913");
        end

        914 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   914");
        end

        915 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   915");
        end

        916 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   916");
        end

        917 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   917");
        end

        918 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   918");
        end

        919 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   919");
        end

        920 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   920");
        end

        921 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   921");
        end

        922 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   922");
        end

        923 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   923");
        end

        924 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   924");
        end

        925 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   925");
        end

        926 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   926");
        end

        927 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   927");
        end

        928 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   928");
        end

        929 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   929");
        end

        930 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   930");
        end

        931 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   931");
        end

        932 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   932");
        end

        933 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   933");
        end

        934 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   934");
        end

        935 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   935");
        end

        936 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   936");
        end

        937 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   937");
        end

        938 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   938");
        end

        939 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   939");
        end

        940 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   940");
        end

        941 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   941");
        end

        942 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   942");
        end

        943 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   943");
        end

        944 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   944");
        end

        945 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   945");
        end

        946 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   946");
        end

        947 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   947");
        end

        948 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   948");
        end

        949 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   949");
        end

        950 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   950");
        end

        951 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   951");
        end

        952 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   952");
        end

        953 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   953");
        end

        954 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   954");
        end

        955 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   955");
        end

        956 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   956");
        end

        957 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   957");
        end

        958 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   958");
        end

        959 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   959");
        end

        960 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   960");
        end

        961 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   961");
        end

        962 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   962");
        end

        963 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   963");
        end

        964 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   964");
        end

        965 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   965");
        end

        966 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   966");
        end

        967 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   967");
        end

        968 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   968");
        end

        969 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   969");
        end

        970 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   970");
        end

        971 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   971");
        end

        972 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   972");
        end

        973 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   973");
        end

        974 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   974");
        end

        975 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   975");
        end

        976 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   976");
        end

        977 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   977");
        end

        978 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   978");
        end

        979 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   979");
        end

        980 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   980");
        end

        981 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   981");
        end

        982 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   982");
        end

        983 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   983");
        end

        984 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   984");
        end

        985 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   985");
        end

        986 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   986");
        end

        987 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   987");
        end

        988 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   988");
        end

        989 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   989");
        end

        990 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   990");
        end

        991 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   991");
        end

        992 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   992");
        end

        993 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   993");
        end

        994 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   994");
        end

        995 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   995");
        end

        996 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   996");
        end

        997 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   997");
        end

        998 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   998");
        end

        999 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   999");
        end

       1000 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1000");
        end

       1001 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1001");
        end

       1002 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1002");
        end

       1003 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1003");
        end

       1004 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1004");
        end

       1005 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1005");
        end

       1006 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1006");
        end

       1007 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1007");
        end

       1008 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1008");
        end

       1009 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1009");
        end

       1010 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1010");
        end

       1011 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1011");
        end

       1012 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1012");
        end

       1013 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1013");
        end

       1014 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1014");
        end

       1015 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1015");
        end

       1016 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1016");
        end

       1017 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1017");
        end

       1018 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1018");
        end

       1019 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1019");
        end

       1020 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1020");
        end

       1021 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1021");
        end

       1022 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1022");
        end

       1023 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1023");
        end

       1024 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1024");
        end

       1025 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1025");
        end

       1026 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1026");
        end

       1027 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1027");
        end

       1028 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1028");
        end

       1029 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1029");
        end

       1030 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1030");
        end

       1031 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1031");
        end

       1032 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1032");
        end

       1033 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1033");
        end

       1034 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1034");
        end

       1035 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1035");
        end

       1036 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1036");
        end

       1037 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1037");
        end

       1038 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1038");
        end

       1039 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1039");
        end

       1040 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1040");
        end

       1041 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1041");
        end

       1042 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1042");
        end

       1043 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1043");
        end

       1044 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1044");
        end

       1045 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1045");
        end

       1046 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1046");
        end

       1047 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1047");
        end

       1048 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1048");
        end

       1049 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1049");
        end

       1050 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1050");
        end

       1051 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1051");
        end

       1052 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1052");
        end

       1053 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1053");
        end

       1054 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1054");
        end

       1055 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1055");
        end

       1056 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1056");
        end

       1057 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1057");
        end

       1058 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1058");
        end

       1059 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1059");
        end

       1060 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1060");
        end

       1061 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1061");
        end

       1062 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1062");
        end

       1063 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1063");
        end

       1064 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1064");
        end

       1065 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1065");
        end

       1066 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1066");
        end

       1067 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1067");
        end

       1068 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1068");
        end

       1069 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1069");
        end

       1070 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1070");
        end

       1071 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1071");
        end

       1072 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1072");
        end

       1073 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1073");
        end

       1074 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1074");
        end

       1075 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1075");
        end

       1076 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1076");
        end

       1077 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1077");
        end

       1078 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1078");
        end

       1079 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1079");
        end

       1080 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1080");
        end

       1081 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1081");
        end

       1082 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1082");
        end

       1083 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1083");
        end

       1084 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1084");
        end

       1085 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1085");
        end

       1086 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1086");
        end

       1087 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1087");
        end

       1088 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1088");
        end

       1089 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1089");
        end

       1090 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1090");
        end

       1091 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1091");
        end

       1092 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1092");
        end

       1093 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1093");
        end

       1094 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1094");
        end

       1095 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1095");
        end

       1096 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1096");
        end

       1097 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1097");
        end

       1098 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1098");
        end

       1099 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1099");
        end

       1100 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1100");
        end

       1101 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1101");
        end

       1102 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1102");
        end

       1103 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1103");
        end

       1104 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1104");
        end

       1105 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1105");
        end

       1106 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1106");
        end

       1107 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1107");
        end

       1108 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1108");
        end

       1109 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1109");
        end

       1110 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1110");
        end

       1111 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1111");
        end

       1112 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1112");
        end

       1113 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1113");
        end

       1114 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1114");
        end

       1115 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1115");
        end

       1116 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1116");
        end

       1117 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1117");
        end

       1118 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1118");
        end

       1119 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1119");
        end

       1120 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1120");
        end

       1121 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1121");
        end

       1122 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1122");
        end

       1123 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1123");
        end

       1124 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1124");
        end

       1125 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1125");
        end

       1126 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1126");
        end

       1127 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1127");
        end

       1128 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1128");
        end

       1129 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1129");
        end

       1130 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1130");
        end

       1131 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1131");
        end

       1132 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1132");
        end

       1133 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1133");
        end

       1134 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1134");
        end

       1135 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1135");
        end

       1136 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1136");
        end

       1137 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1137");
        end

       1138 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1138");
        end

       1139 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1139");
        end

       1140 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1140");
        end

       1141 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1141");
        end

       1142 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1142");
        end

       1143 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1143");
        end

       1144 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1144");
        end

       1145 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1145");
        end

       1146 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1146");
        end

       1147 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1147");
        end

       1148 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1148");
        end

       1149 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1149");
        end

       1150 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
          // $display("Should not be executed  1150");
        end

       1151 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1151");
        end

       1152 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1152");
        end

       1153 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1153");
        end

       1154 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1154");
        end

       1155 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1155");
        end

       1156 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1156");
        end

       1157 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1157");
        end

       1158 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1158");
        end

       1159 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1159");
        end

       1160 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1160");
        end

       1161 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1161");
        end

       1162 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1162");
        end

       1163 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1163");
        end

       1164 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1164");
        end

       1165 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1165");
        end

       1166 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1166");
        end

       1167 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1167");
        end

       1168 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1168");
        end

       1169 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1169");
        end

       1170 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1170");
        end

       1171 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1171");
        end

       1172 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1172");
        end

       1173 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1173");
        end

       1174 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1174");
        end

       1175 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1175");
        end

       1176 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1176");
        end

       1177 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1177");
        end

       1178 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1178");
        end

       1179 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1179");
        end

       1180 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
          // $display("Should not be executed  1180");
        end

       1181 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1181");
        end

       1182 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
          // $display("Should not be executed  1182");
        end

       1183 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1183");
        end

       1184 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1184");
        end

       1185 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1185");
        end

       1186 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1186");
        end

       1187 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1187");
        end

       1188 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1188");
        end

       1189 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1189");
        end

       1190 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1190");
        end

       1191 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1191");
        end

       1192 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1192");
        end

       1193 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1193");
        end

       1194 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1194");
        end

       1195 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1195");
        end

       1196 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1196");
        end

       1197 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1197");
        end

       1198 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1198");
        end

       1199 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1199");
        end

       1200 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1200");
        end

       1201 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1201");
        end

       1202 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1202");
        end

       1203 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1203");
        end

       1204 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1204");
        end

       1205 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1205");
        end

       1206 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1206");
        end

       1207 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1207");
        end

       1208 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1208");
        end

       1209 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1209");
        end

       1210 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1210");
        end

       1211 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1211");
        end

       1212 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1212");
        end

       1213 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1213");
        end

       1214 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1214");
        end

       1215 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1215");
        end

       1216 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1216");
        end

       1217 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1217");
        end

       1218 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1218");
        end

       1219 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1219");
        end

       1220 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1220");
        end

       1221 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1221");
        end

       1222 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1222");
        end

       1223 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1223");
        end

       1224 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1224");
        end

       1225 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1225");
        end

       1226 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1226");
        end

       1227 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1227");
        end

       1228 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1228");
        end

       1229 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1229");
        end

       1230 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1230");
        end

       1231 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1231");
        end

       1232 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1232");
        end

       1233 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1233");
        end

       1234 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1234");
        end

       1235 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1235");
        end

       1236 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1236");
        end

       1237 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1237");
        end

       1238 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1238");
        end

       1239 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1239");
        end

       1240 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1240");
        end

       1241 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1241");
        end

       1242 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1242");
        end

       1243 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1243");
        end

       1244 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1244");
        end

       1245 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1245");
        end

       1246 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1246");
        end

       1247 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1247");
        end

       1248 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1248");
        end

       1249 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1249");
        end

       1250 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1250");
        end

       1251 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1251");
        end

       1252 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1252");
        end

       1253 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1253");
        end

       1254 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1254");
        end

       1255 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1255");
        end

       1256 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1256");
        end

       1257 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1257");
        end

       1258 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1258");
        end

       1259 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1259");
        end

       1260 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1260");
        end

       1261 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1261");
        end

       1262 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1262");
        end

       1263 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1263");
        end

       1264 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1264");
        end

       1265 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1265");
        end

       1266 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1266");
        end

       1267 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1267");
        end

       1268 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1268");
        end

       1269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1269");
        end

       1270 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1270");
        end

       1271 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1271");
        end

       1272 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1272");
        end

       1273 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1273");
        end

       1274 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1274");
        end

       1275 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1275");
        end

       1276 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1276");
        end

       1277 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1277");
        end

       1278 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1278");
        end

       1279 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1279");
        end

       1280 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1280");
        end

       1281 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1281");
        end

       1282 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1282");
        end

       1283 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1283");
        end

       1284 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1284");
        end

       1285 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1285");
        end

       1286 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1286");
        end

       1287 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1287");
        end

       1288 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1288");
        end

       1289 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1289");
        end

       1290 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1290");
        end

       1291 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1291");
        end

       1292 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1292");
        end

       1293 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1293");
        end

       1294 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1294");
        end

       1295 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1295");
        end

       1296 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1296");
        end

       1297 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1297");
        end

       1298 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1298");
        end

       1299 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1299");
        end

       1300 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1300");
        end

       1301 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1301");
        end

       1302 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1302");
        end

       1303 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1303");
        end

       1304 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1304");
        end

       1305 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1305");
        end

       1306 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1306");
        end

       1307 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1307");
        end

       1308 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1308");
        end

       1309 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1309");
        end

       1310 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1310");
        end

       1311 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1311");
        end

       1312 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1312");
        end

       1313 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1313");
        end

       1314 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1314");
        end

       1315 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1315");
        end

       1316 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1316");
        end

       1317 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1317");
        end

       1318 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1318");
        end

       1319 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1319");
        end

       1320 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1320");
        end

       1321 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1321");
        end

       1322 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1322");
        end

       1323 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1323");
        end

       1324 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1324");
        end

       1325 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1325");
        end

       1326 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1326");
        end

       1327 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1327");
        end

       1328 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1328");
        end

       1329 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1329");
        end

       1330 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1330");
        end

       1331 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1331");
        end

       1332 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1332");
        end

       1333 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1333");
        end

       1334 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1334");
        end

       1335 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1335");
        end

       1336 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1336");
        end

       1337 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1337");
        end

       1338 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1338");
        end

       1339 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1339");
        end

       1340 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1340");
        end

       1341 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1341");
        end

       1342 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1342");
        end

       1343 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1343");
        end

       1344 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1344");
        end

       1345 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  1345");
        end

       1346 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1346");
        end

       1347 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1347");
        end

       1348 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1348");
        end

       1349 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1349");
        end

       1350 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1350");
        end

       1351 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1351");
        end

       1352 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1352");
        end

       1353 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1353");
        end

       1354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1354");
        end

       1355 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1355");
        end

       1356 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1356");
        end

       1357 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1357");
        end

       1358 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1358");
        end

       1359 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1359");
        end

       1360 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1360");
        end

       1361 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1361");
        end

       1362 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1362");
        end

       1363 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1363");
        end

       1364 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1364");
        end

       1365 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1365");
        end

       1366 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1366");
        end

       1367 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1367");
        end

       1368 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1368");
        end

       1369 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1369");
        end

       1370 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1370");
        end

       1371 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1371");
        end

       1372 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1372");
        end

       1373 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1373");
        end

       1374 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1374");
        end

       1375 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1375");
        end

       1376 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1376");
        end

       1377 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1377");
        end

       1378 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1378");
        end

       1379 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1379");
        end

       1380 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1380");
        end

       1381 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1381");
        end

       1382 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1382");
        end

       1383 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1383");
        end

       1384 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1384");
        end

       1385 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1385");
        end

       1386 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1386");
        end

       1387 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1387");
        end

       1388 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1388");
        end

       1389 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1389");
        end

       1390 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1390");
        end

       1391 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1391");
        end

       1392 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1392");
        end

       1393 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1393");
        end

       1394 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1394");
        end

       1395 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1395");
        end

       1396 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1396");
        end

       1397 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1397");
        end

       1398 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1398");
        end

       1399 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1399");
        end

       1400 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1400");
        end

       1401 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1401");
        end

       1402 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1402");
        end

       1403 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1403");
        end

       1404 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1404");
        end

       1405 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1405");
        end

       1406 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1406");
        end

       1407 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1407");
        end

       1408 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1408");
        end

       1409 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1409");
        end

       1410 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1410");
        end

       1411 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1411");
        end

       1412 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1412");
        end

       1413 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1413");
        end

       1414 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1414");
        end

       1415 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1415");
        end

       1416 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1416");
        end

       1417 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1417");
        end

       1418 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1418");
        end

       1419 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1419");
        end

       1420 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1420");
        end

       1421 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1421");
        end

       1422 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1422");
        end

       1423 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1423");
        end

       1424 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1424");
        end

       1425 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1425");
        end

       1426 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1426");
        end

       1427 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1427");
        end

       1428 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1428");
        end

       1429 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1429");
        end

       1430 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1430");
        end

       1431 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1431");
        end

       1432 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1432");
        end

       1433 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1433");
        end

       1434 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1434");
        end

       1435 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1435");
        end

       1436 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1436");
        end

       1437 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1437");
        end

       1438 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1438");
        end

       1439 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1439");
        end

       1440 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1440");
        end

       1441 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1441");
        end

       1442 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1442");
        end

       1443 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1443");
        end

       1444 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1444");
        end

       1445 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1445");
        end

       1446 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1446");
        end

       1447 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1447");
        end

       1448 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1448");
        end

       1449 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1449");
        end

       1450 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1450");
        end

       1451 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1451");
        end

       1452 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1452");
        end

       1453 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1453");
        end

       1454 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1454");
        end

       1455 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1455");
        end

       1456 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1456");
        end

       1457 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1457");
        end

       1458 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1458");
        end

       1459 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1459");
        end

       1460 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1460");
        end

       1461 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1461");
        end

       1462 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1462");
        end

       1463 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1463");
        end

       1464 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1464");
        end

       1465 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1465");
        end

       1466 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1466");
        end

       1467 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1467");
        end

       1468 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1468");
        end

       1469 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1469");
        end

       1470 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1470");
        end

       1471 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1471");
        end

       1472 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1472");
        end

       1473 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1473");
        end

       1474 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1474");
        end

       1475 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1475");
        end

       1476 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1476");
        end

       1477 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1477");
        end

       1478 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1478");
        end

       1479 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1479");
        end

       1480 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1480");
        end

       1481 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1481");
        end

       1482 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1482");
        end

       1483 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1483");
        end

       1484 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1484");
        end

       1485 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1485");
        end

       1486 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1486");
        end

       1487 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1487");
        end

       1488 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1488");
        end

       1489 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1489");
        end

       1490 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1490");
        end

       1491 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1491");
        end

       1492 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1492");
        end

       1493 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1493");
        end

       1494 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1494");
        end

       1495 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1495");
        end

       1496 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1496");
        end

       1497 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1497");
        end

       1498 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1498");
        end

       1499 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1499");
        end

       1500 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1500");
        end

       1501 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1501");
        end

       1502 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1502");
        end

       1503 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1503");
        end

       1504 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1504");
        end

       1505 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1505");
        end

       1506 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1506");
        end

       1507 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1507");
        end

       1508 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1508");
        end

       1509 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1509");
        end

       1510 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1510");
        end

       1511 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1511");
        end

       1512 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1512");
        end

       1513 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1513");
        end

       1514 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1514");
        end

       1515 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1515");
        end

       1516 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1516");
        end

       1517 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1517");
        end

       1518 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1518");
        end

       1519 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1519");
        end

       1520 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1520");
        end

       1521 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1521");
        end

       1522 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1522");
        end

       1523 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1523");
        end

       1524 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1524");
        end

       1525 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1525");
        end

       1526 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1526");
        end

       1527 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1527");
        end

       1528 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1528");
        end

       1529 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1529");
        end

       1530 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1530");
        end

       1531 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1531");
        end

       1532 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1532");
        end

       1533 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1533");
        end

       1534 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1534");
        end

       1535 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1535");
        end

       1536 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1536");
        end

       1537 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1537");
        end

       1538 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1538");
        end

       1539 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1539");
        end

       1540 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1540");
        end

       1541 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1541");
        end

       1542 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1542");
        end

       1543 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1543");
        end

       1544 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1544");
        end

       1545 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1545");
        end

       1546 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1546");
        end

       1547 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1547");
        end

       1548 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1548");
        end

       1549 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1549");
        end

       1550 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1550");
        end

       1551 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1551");
        end

       1552 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1552");
        end

       1553 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1553");
        end

       1554 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1554");
        end

       1555 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1555");
        end

       1556 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1556");
        end

       1557 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1557");
        end

       1558 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1558");
        end

       1559 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1559");
        end

       1560 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1560");
        end

       1561 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1561");
        end

       1562 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1562");
        end

       1563 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1563");
        end

       1564 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1564");
        end

       1565 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1565");
        end

       1566 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1566");
        end

       1567 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1567");
        end

       1568 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1568");
        end

       1569 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1569");
        end

       1570 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1570");
        end

       1571 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1571");
        end

       1572 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1572");
        end

       1573 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1573");
        end

       1574 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1574");
        end

       1575 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1575");
        end

       1576 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1576");
        end

       1577 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1577");
        end

       1578 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1578");
        end

       1579 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1579");
        end

       1580 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1580");
        end

       1581 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1581");
        end

       1582 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1582");
        end

       1583 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1583");
        end

       1584 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1584");
        end

       1585 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1585");
        end

       1586 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1586");
        end

       1587 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1587");
        end

       1588 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1588");
        end

       1589 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1589");
        end

       1590 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1590");
        end

       1591 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1591");
        end

       1592 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1592");
        end

       1593 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1593");
        end

       1594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1594");
        end

       1595 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1595");
        end

       1596 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1596");
        end

       1597 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1597");
        end

       1598 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1598");
        end

       1599 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1599");
        end

       1600 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1600");
        end

       1601 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1601");
        end

       1602 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1602");
        end

       1603 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1603");
        end

       1604 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1604");
        end

       1605 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1605");
        end

       1606 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1606");
        end

       1607 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1607");
        end

       1608 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1608");
        end

       1609 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1609");
        end

       1610 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1610");
        end

       1611 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1611");
        end

       1612 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1612");
        end

       1613 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1613");
        end

       1614 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1614");
        end

       1615 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1615");
        end

       1616 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1616");
        end

       1617 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1617");
        end

       1618 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1618");
        end

       1619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1619");
        end

       1620 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1620");
        end

       1621 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1621");
        end

       1622 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1622");
        end

       1623 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1623");
        end

       1624 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1624");
        end

       1625 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1625");
        end

       1626 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1626");
        end

       1627 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1627");
        end

       1628 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1628");
        end

       1629 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1629");
        end

       1630 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1630");
        end

       1631 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1631");
        end

       1632 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1632");
        end

       1633 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1633");
        end

       1634 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1634");
        end

       1635 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1635");
        end

       1636 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1636");
        end

       1637 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1637");
        end

       1638 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1638");
        end

       1639 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1639");
        end

       1640 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1640");
        end

       1641 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1641");
        end

       1642 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1642");
        end

       1643 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1643");
        end

       1644 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1644");
        end

       1645 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1645");
        end

       1646 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1646");
        end

       1647 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1647");
        end

       1648 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1648");
        end

       1649 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1649");
        end

       1650 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  1650");
        end

       1651 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1651");
        end

       1652 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1652");
        end

       1653 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1653");
        end

       1654 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1654");
        end

       1655 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1655");
        end

       1656 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1656");
        end

       1657 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1657");
        end

       1658 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1658");
        end

       1659 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1659");
        end

       1660 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1660");
        end

       1661 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1661");
        end

       1662 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1662");
        end

       1663 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1663");
        end

       1664 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1664");
        end

       1665 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1665");
        end

       1666 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1666");
        end

       1667 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1667");
        end

       1668 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1668");
        end

       1669 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1669");
        end

       1670 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1670");
        end

       1671 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1671");
        end

       1672 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1672");
        end

       1673 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1673");
        end

       1674 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1674");
        end

       1675 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1675");
        end

       1676 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1676");
        end

       1677 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1677");
        end

       1678 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1678");
        end

       1679 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1679");
        end

       1680 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1680");
        end

       1681 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1681");
        end

       1682 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1682");
        end

       1683 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1683");
        end

       1684 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1684");
        end

       1685 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1685");
        end

       1686 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1686");
        end

       1687 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1687");
        end

       1688 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1688");
        end

       1689 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1689");
        end

       1690 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1690");
        end

       1691 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1691");
        end

       1692 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1692");
        end

       1693 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1693");
        end

       1694 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1694");
        end

       1695 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1695");
        end

       1696 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1696");
        end

       1697 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1697");
        end

       1698 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1698");
        end

       1699 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1699");
        end

       1700 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1700");
        end

       1701 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1701");
        end

       1702 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1702");
        end

       1703 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1703");
        end

       1704 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1704");
        end

       1705 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1705");
        end

       1706 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1706");
        end

       1707 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1707");
        end

       1708 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1708");
        end

       1709 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1709");
        end

       1710 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1710");
        end

       1711 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1711");
        end

       1712 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1712");
        end

       1713 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1713");
        end

       1714 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
          // $display("Should not be executed  1714");
        end

       1715 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1715");
        end

       1716 :
        begin                                                                   // shiftRight
          //$display("AAAA %4d %4d shiftRight", steps, ip);
          // $display("Should not be executed  1716");
        end

       1717 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1717");
        end

       1718 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1718");
        end

       1719 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1719");
        end

       1720 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1720");
        end

       1721 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
          // $display("Should not be executed  1721");
        end

       1722 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1722");
        end

       1723 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1723");
        end

       1724 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1724");
        end

       1725 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1725");
        end

       1726 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1726");
        end

       1727 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1727");
        end

       1728 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1728");
        end

       1729 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1729");
        end

       1730 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1730");
        end

       1731 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1731");
        end

       1732 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1732");
        end

       1733 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1733");
        end

       1734 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1734");
        end

       1735 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1735");
        end

       1736 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1736");
        end

       1737 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1737");
        end

       1738 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1738");
        end

       1739 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1739");
        end

       1740 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1740");
        end

       1741 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1741");
        end

       1742 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1742");
        end

       1743 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1743");
        end

       1744 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1744");
        end

       1745 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1745");
        end

       1746 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1746");
        end

       1747 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1747");
        end

       1748 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1748");
        end

       1749 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1749");
        end

       1750 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1750");
        end

       1751 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1751");
        end

       1752 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1752");
        end

       1753 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1753");
        end

       1754 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1754");
        end

       1755 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1755");
        end

       1756 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1756");
        end

       1757 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1757");
        end

       1758 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1758");
        end

       1759 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1759");
        end

       1760 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1760");
        end

       1761 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1761");
        end

       1762 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1762");
        end

       1763 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1763");
        end

       1764 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1764");
        end

       1765 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1765");
        end

       1766 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1766");
        end

       1767 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1767");
        end

       1768 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1768");
        end

       1769 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1769");
        end

       1770 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1770");
        end

       1771 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1771");
        end

       1772 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1772");
        end

       1773 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1773");
        end

       1774 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1774");
        end

       1775 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1775");
        end

       1776 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1776");
        end

       1777 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1777");
        end

       1778 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1778");
        end

       1779 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1779");
        end

       1780 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1780");
        end

       1781 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1781");
        end

       1782 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1782");
        end

       1783 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1783");
        end

       1784 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1784");
        end

       1785 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1785");
        end

       1786 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1786");
        end

       1787 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1787");
        end

       1788 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1788");
        end

       1789 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1789");
        end

       1790 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1790");
        end

       1791 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1791");
        end

       1792 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1792");
        end

       1793 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1793");
        end

       1794 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1794");
        end

       1795 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1795");
        end

       1796 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1796");
        end

       1797 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1797");
        end

       1798 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1798");
        end

       1799 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1799");
        end

       1800 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1800");
        end

       1801 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1801");
        end

       1802 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1802");
        end

       1803 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1803");
        end

       1804 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1804");
        end

       1805 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1805");
        end

       1806 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1806");
        end

       1807 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1807");
        end

       1808 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1808");
        end

       1809 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1809");
        end

       1810 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1810");
        end

       1811 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1811");
        end

       1812 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1812");
        end

       1813 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1813");
        end

       1814 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1814");
        end

       1815 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1815");
        end

       1816 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1816");
        end

       1817 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1817");
        end

       1818 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1818");
        end

       1819 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1819");
        end

       1820 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1820");
        end

       1821 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1821");
        end

       1822 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1822");
        end

       1823 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1823");
        end

       1824 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1824");
        end

       1825 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1825");
        end

       1826 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1826");
        end

       1827 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1827");
        end

       1828 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1828");
        end

       1829 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1829");
        end

       1830 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1830");
        end

       1831 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1831");
        end

       1832 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1832");
        end

       1833 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1833");
        end

       1834 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1834");
        end

       1835 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1835");
        end

       1836 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1836");
        end

       1837 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1837");
        end

       1838 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1838");
        end

       1839 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1839");
        end

       1840 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1840");
        end

       1841 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1841");
        end

       1842 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1842");
        end

       1843 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1843");
        end

       1844 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1844");
        end

       1845 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1845");
        end

       1846 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1846");
        end

       1847 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1847");
        end

       1848 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1848");
        end

       1849 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1849");
        end

       1850 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1850");
        end

       1851 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1851");
        end

       1852 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1852");
        end

       1853 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1853");
        end

       1854 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1854");
        end

       1855 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1855");
        end

       1856 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1856");
        end

       1857 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1857");
        end

       1858 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1858");
        end

       1859 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1859");
        end

       1860 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1860");
        end

       1861 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1861");
        end

       1862 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1862");
        end

       1863 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1863");
        end

       1864 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1864");
        end

       1865 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1865");
        end

       1866 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1866");
        end

       1867 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1867");
        end

       1868 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1868");
        end

       1869 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1869");
        end

       1870 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1870");
        end

       1871 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1871");
        end

       1872 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1872");
        end

       1873 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1873");
        end

       1874 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1874");
        end

       1875 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1875");
        end

       1876 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1876");
        end

       1877 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1877");
        end

       1878 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1878");
        end

       1879 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed  1879");
        end

       1880 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1880");
        end

       1881 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1881");
        end

       1882 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1882");
        end

       1883 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed  1883");
        end

       1884 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1884");
        end

       1885 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1885");
        end

       1886 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1886");
        end

       1887 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1887");
        end

       1888 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1888");
        end

       1889 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1889");
        end

       1890 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1890");
        end

       1891 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1891");
        end

       1892 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1892");
        end

       1893 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1893");
        end

       1894 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1894");
        end

       1895 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1895");
        end

       1896 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1896");
        end

       1897 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1897");
        end

       1898 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1898");
        end

       1899 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1899");
        end

       1900 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1900");
        end

       1901 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1901");
        end

       1902 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1902");
        end

       1903 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1903");
        end

       1904 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1904");
        end

       1905 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1905");
        end

       1906 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1906");
        end

       1907 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1907");
        end

       1908 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1908");
        end

       1909 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1909");
        end

       1910 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1910");
        end

       1911 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1911");
        end

       1912 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1912");
        end

       1913 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1913");
        end

       1914 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1914");
        end

       1915 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1915");
        end

       1916 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1916");
        end

       1917 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1917");
        end

       1918 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed  1918");
        end

       1919 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1919");
        end

       1920 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1920");
        end

       1921 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1921");
        end

       1922 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1922");
        end

       1923 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1923");
        end

       1924 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1924");
        end

       1925 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1925");
        end

       1926 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1926");
        end

       1927 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1927");
        end

       1928 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1928");
        end

       1929 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1929");
        end

       1930 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1930");
        end

       1931 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1931");
        end

       1932 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1932");
        end

       1933 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1933");
        end

       1934 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1934");
        end

       1935 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1935");
        end

       1936 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1936");
        end

       1937 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1937");
        end

       1938 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1938");
        end

       1939 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1939");
        end

       1940 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1940");
        end

       1941 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1941");
        end

       1942 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1942");
        end

       1943 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1943");
        end

       1944 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1944");
        end

       1945 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1945");
        end

       1946 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1946");
        end

       1947 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1947");
        end

       1948 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1948");
        end

       1949 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1949");
        end

       1950 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1950");
        end

       1951 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1951");
        end

       1952 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1952");
        end

       1953 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1953");
        end

       1954 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1954");
        end

       1955 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1955");
        end

       1956 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1956");
        end

       1957 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1957");
        end

       1958 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1958");
        end

       1959 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1959");
        end

       1960 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1960");
        end

       1961 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1961");
        end

       1962 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1962");
        end

       1963 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1963");
        end

       1964 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1964");
        end

       1965 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1965");
        end

       1966 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1966");
        end

       1967 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1967");
        end

       1968 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1968");
        end

       1969 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1969");
        end

       1970 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1970");
        end

       1971 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1971");
        end

       1972 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1972");
        end

       1973 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1973");
        end

       1974 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1974");
        end

       1975 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1975");
        end

       1976 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1976");
        end

       1977 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1977");
        end

       1978 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1978");
        end

       1979 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1979");
        end

       1980 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1980");
        end

       1981 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1981");
        end

       1982 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1982");
        end

       1983 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1983");
        end

       1984 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1984");
        end

       1985 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1985");
        end

       1986 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1986");
        end

       1987 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1987");
        end

       1988 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1988");
        end

       1989 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1989");
        end

       1990 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1990");
        end

       1991 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1991");
        end

       1992 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1992");
        end

       1993 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1993");
        end

       1994 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1994");
        end

       1995 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1995");
        end

       1996 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1996");
        end

       1997 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1997");
        end

       1998 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1998");
        end

       1999 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1999");
        end

       2000 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2000");
        end

       2001 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2001");
        end

       2002 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2002");
        end

       2003 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2003");
        end

       2004 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2004");
        end

       2005 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2005");
        end

       2006 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2006");
        end

       2007 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2007");
        end

       2008 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2008");
        end

       2009 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2009");
        end

       2010 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2010");
        end

       2011 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2011");
        end

       2012 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2012");
        end

       2013 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2013");
        end

       2014 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2014");
        end

       2015 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2015");
        end

       2016 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2016");
        end

       2017 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2017");
        end

       2018 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2018");
        end

       2019 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2019");
        end

       2020 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2020");
        end

       2021 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2021");
        end

       2022 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2022");
        end

       2023 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2023");
        end

       2024 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2024");
        end

       2025 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2025");
        end

       2026 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2026");
        end

       2027 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2027");
        end

       2028 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2028");
        end

       2029 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2029");
        end

       2030 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2030");
        end

       2031 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2031");
        end

       2032 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2032");
        end

       2033 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2033");
        end

       2034 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2034");
        end

       2035 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2035");
        end

       2036 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2036");
        end

       2037 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2037");
        end

       2038 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2038");
        end

       2039 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2039");
        end

       2040 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2040");
        end

       2041 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2041");
        end

       2042 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2042");
        end

       2043 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2043");
        end

       2044 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2044");
        end

       2045 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2045");
        end

       2046 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2046");
        end

       2047 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2047");
        end

       2048 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2048");
        end

       2049 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2049");
        end

       2050 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2050");
        end

       2051 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2051");
        end

       2052 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2052");
        end

       2053 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2053");
        end

       2054 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2054");
        end

       2055 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2055");
        end

       2056 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2056");
        end

       2057 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2057");
        end

       2058 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2058");
        end

       2059 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2059");
        end

       2060 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2060");
        end

       2061 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2061");
        end

       2062 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2062");
        end

       2063 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2063");
        end

       2064 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2064");
        end

       2065 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2065");
        end

       2066 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2066");
        end

       2067 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2067");
        end

       2068 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2068");
        end

       2069 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2069");
        end

       2070 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2070");
        end

       2071 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2071");
        end

       2072 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2072");
        end

       2073 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2073");
        end

       2074 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2074");
        end

       2075 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2075");
        end

       2076 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2076");
        end

       2077 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2077");
        end

       2078 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2078");
        end

       2079 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2079");
        end

       2080 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2080");
        end

       2081 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2081");
        end

       2082 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2082");
        end

       2083 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2083");
        end

       2084 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2084");
        end

       2085 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2085");
        end

       2086 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2086");
        end

       2087 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2087");
        end

       2088 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2088");
        end

       2089 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2089");
        end

       2090 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2090");
        end

       2091 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2091");
        end

       2092 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2092");
        end

       2093 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2093");
        end

       2094 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2094");
        end

       2095 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2095");
        end

       2096 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2096");
        end

       2097 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2097");
        end

       2098 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2098");
        end

       2099 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2099");
        end

       2100 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2100");
        end

       2101 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2101");
        end

       2102 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2102");
        end

       2103 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2103");
        end

       2104 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2104");
        end

       2105 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2105");
        end

       2106 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2106");
        end

       2107 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2107");
        end

       2108 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2108");
        end

       2109 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2109");
        end

       2110 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2110");
        end

       2111 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2111");
        end

       2112 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2112");
        end

       2113 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2113");
        end

       2114 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2114");
        end

       2115 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2115");
        end

       2116 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2116");
        end

       2117 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2117");
        end

       2118 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2118");
        end

       2119 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2119");
        end

       2120 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2120");
        end

       2121 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2121");
        end

       2122 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2122");
        end

       2123 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2123");
        end

       2124 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2124");
        end

       2125 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2125");
        end

       2126 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2126");
        end

       2127 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2127");
        end

       2128 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2128");
        end

       2129 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2129");
        end

       2130 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2130");
        end

       2131 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2131");
        end

       2132 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2132");
        end

       2133 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2133");
        end

       2134 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2134");
        end

       2135 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2135");
        end

       2136 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2136");
        end

       2137 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2137");
        end

       2138 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2138");
        end

       2139 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2139");
        end

       2140 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2140");
        end

       2141 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2141");
        end

       2142 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2142");
        end

       2143 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2143");
        end

       2144 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2144");
        end

       2145 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2145");
        end

       2146 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2146");
        end

       2147 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2147");
        end

       2148 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2148");
        end

       2149 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2149");
        end

       2150 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2150");
        end

       2151 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2151");
        end

       2152 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2152");
        end

       2153 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2153");
        end

       2154 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2154");
        end

       2155 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2155");
        end

       2156 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2156");
        end

       2157 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2157");
        end

       2158 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2158");
        end

       2159 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2159");
        end

       2160 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2160");
        end

       2161 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2161");
        end

       2162 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2162");
        end

       2163 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2163");
        end

       2164 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2164");
        end

       2165 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2165");
        end

       2166 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2166");
        end

       2167 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2167");
        end

       2168 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2168");
        end

       2169 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2169");
        end

       2170 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2170");
        end

       2171 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2171");
        end

       2172 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2172");
        end

       2173 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2173");
        end

       2174 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2174");
        end

       2175 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2175");
        end

       2176 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2176");
        end

       2177 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2177");
        end

       2178 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2178");
        end

       2179 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2180;
        end

       2180 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[1];
              ip = 2181;
              heapClock = ~ heapClock;
        end
      endcase
      success  = 1;
      finished = steps >     73;
    end
  end

endmodule
