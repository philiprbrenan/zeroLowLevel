// Check double frees, over allocation
// Check access to unallocated arrays or elements
// Check push overflow, pop underflow
// Next Message 10000280
`define Reset        1  /* Zero all memory sizes                               */
`define Write        2  /* Write an element                                    */
`define Read         3  /* Read an element                                     */
`define Size         4  /* Size of array                                       */
`define Inc          5  /* Increment size of array if possible                 */
`define Dec          6  /* Decrement size of array if possible                 */
`define Index        7  /* Index of element in array                           */
`define Less         8  /* Elements of array less than in                      */
`define Greater      9  /* Elements of array greater than in                   */
`define Up          10  /* Move array up                                       */
`define Down        11  /* Move array down                                     */
`define Long1       12  /* Move long first step                                */
`define Long2       13  /* Move long last  step                                */
`define Push        14  /* Push if possible                                    */
`define Pop         15  /* Pop if possible                                     */
`define Dump        16  /* Dump                                                */
`define Resize      17  /* Resize an array                                     */
`define Alloc       18  /* Allocate a new array before using it                */
`define Free        19  /* Free an array for reuse                             */
`define Add         20  /* Add to an element returning the new value           */
`define AddAfter    21  /* Add to an element returning the previous value      */
`define Subtract    22  /* Subtract to an element returning the new value      */
`define SubAfter    23  /* Subtract to an element returning the previous value */
`define ShiftLeft   24  /* Shift left                                          */
`define ShiftRight  25  /* Shift right                                         */
`define NotLogical  26  /* Not - logical                                       */
`define Not         27  /* Not - bitwise                                       */
`define Or          28  /* Or                                                  */
`define Xor         29  /* Xor                                                 */
`define And         30  /* And                                                 */

module Memory
#(parameter integer ADDRESS_BITS =  8,                                          // Number of bits in an address
  parameter integer INDEX_BITS   =  3,                                          // Bits in in an index
  parameter integer DATA_BITS    = 16)                                          // Width of an element in bits
 (input wire                    clock,                                          // Clock to drive array operations
  input wire[7:0]               action,                                         // Operation to be performed on array
  input wire [ADDRESS_BITS-1:0] array,                                          // The number of the array to work on
  input wire [INDEX_BITS  -1:0] index,                                          // Index within array
  input wire [DATA_BITS   -1:0] in,                                             // Input data
  output reg [DATA_BITS   -1:0] out,                                            // Output data
  output reg [31:0]             error);                                         // Error

  parameter integer ARRAY_LENGTH = 2**INDEX_BITS;                               // Maximum index
  parameter integer ARRAYS       = 2**ADDRESS_BITS;                             // Number of memory elements for both arrays and elements

  reg [DATA_BITS   -1:0] memory     [ARRAYS-1:0][ARRAY_LENGTH-1:0];             // Memory containing arrays in fixed blocks
  reg [DATA_BITS   -1:0] copy                   [ARRAY_LENGTH-1:0];             // Copy of one array
  reg [INDEX_BITS    :0] arraySizes [ARRAYS-1:0];                               // Current size of each array
  reg [ADDRESS_BITS-1:0] freedArrays[ARRAYS-1:0];                               // Currently freed arrays
  reg                    allocations[ARRAYS-1:0];                               // Currently allocated arrays

  integer allocatedArrays;                                                      // Arrays allocated
  integer freedArraysTop;                                                       // Top of the freed arrays stack
  integer result;                                                               // Result of each array operation
  integer size;                                                                 // Size of current array
  integer moveLongStartArray;                                                   // Source array of move long
  integer moveLongStartIndex;                                                   // Source index of move long
  integer i, a, b;                                                              // Index

  task checkWriteable(input integer err);                                       // Check a memory is writable
    begin
       error = 0;
       if (array >= allocatedArrays) begin
         //$display("Array has not been allocated, array %d", array);
         error = err;
       end
       if (!allocations[array]) begin
         //$display("Array has been freed, array %d", array);
         error = err + 1;
       end
    end
  endtask

  task checkReadable(input integer err);                                        // Check a memory locationis readable
    begin
       checkWriteable(err);
       if (index >= arraySizes[array]) begin
         //$display("Access outside array bounds, array %d, size: %d, access: %d", array, arraySizes[array], index);
         error = err + 2;
       end
    end
  endtask

  task dump;                                                                    // Dump some memory
    begin
      //$display("    %2d %2d %2d", arraySizes[0], arraySizes[1], arraySizes[2]);
      for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
        //$display("%2d  %2d %2d %2d", i, memory[0][i], memory[1][i], memory[2][i]);
      end
      //$display("    %2d %2d %2d", allocations[0], allocations[1], allocations[2]);
    end
  endtask

  always @(clock) begin                                                             // Each transition
    case(action)                                                                // Decode request
      `Reset: begin                                                             // Reset
        freedArraysTop = 0;                                                     // Free all arrays
        allocatedArrays = 0;
      end

      `Write: begin                                                             // Write
        checkWriteable(10000010);
        if (!error) begin
          memory[array][index] = in;
          if (index >= arraySizes[array] && index < ARRAY_LENGTH) begin
            arraySizes[array] = index + 1;
          end
          out = in;
        end
      end

      `Read: begin                                                              // Read
        checkReadable(10000020);
        if (!error) begin
          out = memory[array][index];
        end
      end

      `Size: begin                                                              // Size
        checkWriteable(10000030);
        if (!error) begin
          out = arraySizes[array];
        end
      end

      `Dec: begin                                                               // Decrement
        checkWriteable(10000040);
        if (!error) begin
          if (arraySizes[array] > 0) arraySizes[array] = arraySizes[array] - 1;
          else begin
            //$display("Attempt to decrement empty array, array %d", array); error = 10000044;
          end
        end
      end

      `Inc: begin                                                               // Increment
        checkWriteable(10000050);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;
          else begin
            //$display("Attempt to decrement full array, array %d", array);  error = 10000054;
          end
        end
      end

      `Index: begin                                                             // Index
        checkWriteable(10000060);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] == in) result = i + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Less: begin                                                              // Count less
        checkWriteable(10000070);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] < in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Greater: begin                                                           // Count greater
        checkWriteable(10000080);
        if (!error) begin
          result = 0;
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin
            if (i < size && memory[array][i] > in) result = result + 1;
////$display("AAAA %d %d %d %d %d", i, size, memory[array][i], in, result);
          end
          out = result;
        end
      end

      `Down: begin                                                              // Down
        checkWriteable(10000270);
        if (!error) begin
          size   = arraySizes[array];
          if (size > 0) begin
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i]; // Copy source array
            for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                       // Move original array up
              if (i > index && i <= size) begin
                memory[array][i-1] = copy[i];
              end
            end
            out = copy[index];                                                  // Return replaced value
            arraySizes[array] = arraySizes[array] - 1;                          // Decrease array size
          end
          else error = 100000274;                                               // Orignal array was emoty so we cannot shift it down
        end
      end

      `Up: begin                                                                // Up
        checkWriteable(10000090);
        if (!error) begin
          size   = arraySizes[array];
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) copy[i] = memory[array][i];   // Copy source array
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Move original array up
            if (i > index && i <= size) begin
              memory[array][i] = copy[i-1];
            end
          end
          memory[array][index] = in;                                            // Insert new value
          if (size < ARRAY_LENGTH) arraySizes[array] = arraySizes[array] + 1;   // Increase array size
        end
      end

      `Long1: begin                                                             // Move long start
        checkReadable(10000100);
        if (!error) begin
          moveLongStartArray = array;                                           // Record source
          moveLongStartIndex = index;
        end
      end

      `Long2: begin                                                             // Move long finish
        checkWriteable(10000110);
        if (!error) begin
          for(i = 0; i < ARRAY_LENGTH; i = i + 1) begin                         // Copy from source to target
            if (i < in && index + i < ARRAY_LENGTH && moveLongStartIndex+i < ARRAY_LENGTH) begin
              memory[array][index+i] = memory[moveLongStartArray][moveLongStartIndex+i];
              if (index+i >= arraySizes[array]) arraySizes[array] = index+i+1;
            end
          end
        end
      end

      `Push: begin                                                              // Push
        checkWriteable(10000120);
        if (!error) begin
          if (arraySizes[array] < ARRAY_LENGTH) begin
            memory[array][arraySizes[array]] = in;
            arraySizes[array] = arraySizes[array] + 1;
          end
          else begin
            //$display("Attempt to push to full array, array %d, value %d", array, in);  error = 10000124;
          end
        end
      end

      `Pop: begin                                                               // Pop
        checkWriteable(10000130);
        if (!error) begin
          if (arraySizes[array] > 0) begin
            arraySizes[array] = arraySizes[array] - 1;
            out = memory[array][arraySizes[array]];
          end
          else begin
            //$display("Attempt to pop empty array, array %d", array); error = 10000134;
          end
        end
      end

      `Dump: begin                                                              // Dump
        dump();
      end

      `Resize: begin                                                            // Resize
        checkWriteable(10000140);
        if (!error) begin
          if (in <= ARRAY_LENGTH) arraySizes[array] = in;
          else begin
            //$display("Attempt to make an array too large, array %d, max %d, size %d", array, ARRAY_LENGTH, in); error = 10000144;
          end
        end
      end

      `Alloc: begin                                                             // Allocate an array
        if (freedArraysTop > 0) begin                                           // Reuse a freed array
          freedArraysTop = freedArraysTop - 1;
          result = freedArrays[freedArraysTop];
        end
        else if (allocatedArrays < ARRAYS-1) begin                              // Allocate a new array - assumes enough memory
          result          = allocatedArrays;
          allocatedArrays = allocatedArrays + 1;
        end
        else begin
          //$display("Out of memory, cannot allocate a new array"); error = 10000270;
        end
        allocations[result] = 1;                                                // Allocated
        arraySizes[result] = 0;                                                 // Empty array
        out = result;
      end

      `Free: begin                                                              // Free an array
        checkWriteable(10000150);
        if (!error) begin
          freedArrays[freedArraysTop] = array;                                  // Relies on the user not re freeing a freed array - we should probably hve another array to prevent this
          allocations[array]          = 0;                                      // No longer allocated
          freedArraysTop = freedArraysTop + 1;
        end
      end

      `Add: begin                                                               // Add to an element
        checkReadable(10000160);
        if (!error) begin
          memory[array][index] = memory[array][index] + in;
          out = memory[array][index];
        end
      end

      `AddAfter: begin                                                          // Add to an element after putting the content of the element on out
        checkReadable(10000170);
        if (!error) begin
        out = memory[array][index];
        memory[array][index] = memory[array][index] + in;
        end
      end

      `Subtract: begin                                                          // Subtract from an element
        checkReadable(10000180);
        if (!error) begin
          memory[array][index] = memory[array][index] - in;
          out = memory[array][index];
        end
      end

      `SubAfter: begin                                                          // Subtract from an element after putting the content of the element on out
        checkReadable(10000190);
        if (!error) begin
          out = memory[array][index];
          memory[array][index] = memory[array][index] - in;
        end
      end

      `ShiftLeft: begin                                                         // Shift left
        checkReadable(10000200);
        if (!error) begin
          memory[array][index] = memory[array][index] << in;
          out = memory[array][index];
        end
      end

      `ShiftRight: begin                                                        // Shift right
        checkReadable(10000210);
        if (!error) begin
          memory[array][index] = memory[array][index] >> in;
          out = memory[array][index];
        end
      end

      `NotLogical: begin                                                        // Not logical
        checkReadable(10000220);
        if (!error) begin
          memory[array][index] = !memory[array][index];
          out = memory[array][index];
        end
      end

      `Not: begin                                                               // Not
        checkReadable(10000230);
        if (!error) begin
          memory[array][index] = ~memory[array][index];
          out = memory[array][index];
        end
      end

      `Or: begin                                                                // Or
        checkReadable(10000240);
        if (!error) begin
          memory[array][index] = memory[array][index] | in;
          out = memory[array][index];
        end
      end

      `Xor: begin                                                               // Xor
        checkReadable(10000250);
        if (!error) begin
          memory[array][index] = memory[array][index] ^ in;
          out = memory[array][index];
        end
      end

      `And: begin                                                               // And
        checkReadable(10000260);
        if (!error) begin
          memory[array][index] = memory[array][index] & in;
          out = memory[array][index];
        end
      end
    endcase
  end
endmodule
//-----------------------------------------------------------------------------
// Fpga test
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga                                                                     // Run test programs
 (input  wire clock,                                                            // Driving clock
  input  wire reset,                                                            // Restart program
  output reg  finished,                                                         // Goes high when the program has finished
  output reg  success);                                                         // Goes high on finish if all the tests passed

  reg                heapClock;                                                 // Clock to drive array operations
  reg [7:0]          heapAction;                                                // Operation to be performed on array
  reg [       8-1:0] heapArray;                                         // The number of the array to work on
  reg [       3-1:0] heapIndex;                                         // Index within array
  reg [      12-1:0] heapIn;                                            // Input data
  reg [      12-1:0] heapOut;                                           // Output data
  reg [31        :0] heapError;                                                 // Error on heap operation if not zero

  Memory                                                                        // Memory module
   #(       8,        3,       12)                          // Address bits, index bits, data bits
    heap(                                                                       // Create heap memory
    .clock  (heapClock),
    .action (heapAction),
    .array  (heapArray),
    .index  (heapIndex),
    .in     (heapIn),
    .out    (heapOut),
    .error  (heapError)
  );
  parameter integer NIn =      107;                                           // Size of input area
  reg [      12-1:0] localMem[    1251-1:0];                       // Local memory
  reg [      12-1:0]   outMem[     107  -1:0];                       // Out channel
  reg [      12-1:0]    inMem[     107   -1:0];                       // In channel

  integer inMemPos;                                                             // Current position in input channel
  integer outMemPos;                                                            // Position in output channel

  integer ip;                                                                   // Instruction pointer
  integer steps;                                                                // Number of steps executed so far
  integer i, j, k;                                                              // A useful counter

  always @(posedge clock, negedge clock) begin                                  // Each instruction
    if (reset) begin
      ip             = 0;
      steps          = 0;
      inMemPos       = 0;
      outMemPos      = 0;
      finished       = 0;
      success        = 0;

      inMem[0] = 72;
      inMem[1] = 103;
      inMem[2] = 3;
      inMem[3] = 89;
      inMem[4] = 49;
      inMem[5] = 6;
      inMem[6] = 38;
      inMem[7] = 91;
      inMem[8] = 21;
      inMem[9] = 39;
      inMem[10] = 52;
      inMem[11] = 62;
      inMem[12] = 19;
      inMem[13] = 83;
      inMem[14] = 7;
      inMem[15] = 70;
      inMem[16] = 73;
      inMem[17] = 18;
      inMem[18] = 40;
      inMem[19] = 67;
      inMem[20] = 59;
      inMem[21] = 10;
      inMem[22] = 20;
      inMem[23] = 56;
      inMem[24] = 86;
      inMem[25] = 90;
      inMem[26] = 27;
      inMem[27] = 98;
      inMem[28] = 45;
      inMem[29] = 15;
      inMem[30] = 1;
      inMem[31] = 48;
      inMem[32] = 33;
      inMem[33] = 4;
      inMem[34] = 28;
      inMem[35] = 87;
      inMem[36] = 24;
      inMem[37] = 66;
      inMem[38] = 84;
      inMem[39] = 80;
      inMem[40] = 65;
      inMem[41] = 75;
      inMem[42] = 97;
      inMem[43] = 85;
      inMem[44] = 63;
      inMem[45] = 54;
      inMem[46] = 12;
      inMem[47] = 101;
      inMem[48] = 31;
      inMem[49] = 41;
      inMem[50] = 30;
      inMem[51] = 106;
      inMem[52] = 26;
      inMem[53] = 68;
      inMem[54] = 60;
      inMem[55] = 95;
      inMem[56] = 35;
      inMem[57] = 76;
      inMem[58] = 96;
      inMem[59] = 61;
      inMem[60] = 105;
      inMem[61] = 32;
      inMem[62] = 42;
      inMem[63] = 37;
      inMem[64] = 43;
      inMem[65] = 57;
      inMem[66] = 102;
      inMem[67] = 93;
      inMem[68] = 29;
      inMem[69] = 78;
      inMem[70] = 55;
      inMem[71] = 82;
      inMem[72] = 23;
      inMem[73] = 22;
      inMem[74] = 44;
      inMem[75] = 9;
      inMem[76] = 81;
      inMem[77] = 5;
      inMem[78] = 79;
      inMem[79] = 14;
      inMem[80] = 13;
      inMem[81] = 51;
      inMem[82] = 88;
      inMem[83] = 74;
      inMem[84] = 94;
      inMem[85] = 17;
      inMem[86] = 16;
      inMem[87] = 2;
      inMem[88] = 47;
      inMem[89] = 36;
      inMem[90] = 8;
      inMem[91] = 100;
      inMem[92] = 53;
      inMem[93] = 25;
      inMem[94] = 34;
      inMem[95] = 64;
      inMem[96] = 77;
      inMem[97] = 46;
      inMem[98] = 99;
      inMem[99] = 11;
      inMem[100] = 50;
      inMem[101] = 69;
      inMem[102] = 58;
      inMem[103] = 104;
      inMem[104] = 71;
      inMem[105] = 92;
      inMem[106] = 107;
    end
    else begin
      case(ip)

          0 :
        begin                                                                   // start
          //$display("AAAA %4d %4d start", steps, ip);
              heapClock = 0;                                                    // Ready for next operation
              ip = 1;
        end

          1 :
        begin                                                                   // start2
          //$display("AAAA %4d %4d start2", steps, ip);
              heapAction = `Reset;                                          // Ready for next operation
              ip = 2;
              heapClock = ~ heapClock;
        end

          2 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 3;
              heapClock = ~ heapClock;
        end

          3 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[0] = heapOut;
              ip = 4;
        end

          4 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[540] = 3;
              ip = 5;
        end

          5 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[540];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 6;
              heapClock = ~ heapClock;
        end

          6 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[541] = 0;
              ip = 7;
        end

          7 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[541];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 8;
              heapClock = ~ heapClock;
        end

          8 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[542] = 0;
              ip = 9;
        end

          9 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[542];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 10;
              heapClock = ~ heapClock;
        end

         10 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[543] = 0;
              ip = 11;
        end

         11 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[543];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 12;
              heapClock = ~ heapClock;
        end

         12 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 13;
              heapClock = ~ heapClock;
        end

         13 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[1] = heapOut;
              ip = 14;
        end

         14 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 15;
        end

         15 :
        begin                                                                   // inSize
          //$display("AAAA %4d %4d inSize", steps, ip);
              localMem[2] = 107 - inMemPos;
              ip = 16;
        end

         16 :
        begin                                                                   // jFalse
          //$display("AAAA %4d %4d jFalse", steps, ip);
              ip = localMem[2] == 0 ? 2168 : 17;
        end

         17 :
        begin                                                                   // in
          //$display("AAAA %4d %4d in", steps, ip);
              if (inMemPos < 107) begin
                localMem[3] = inMem[inMemPos];
                inMemPos = inMemPos + 1;
              end
              ip = 18;
        end

         18 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 19;
              heapClock = ~ heapClock;
        end

         19 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[544] = heapOut;                                                     // Data retrieved from heap memory
              ip = 20;
              heapClock = ~ heapClock;
        end

         20 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[4] = localMem[544];
              ip = 21;
        end

         21 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[5] = localMem[3] + localMem[3];
              ip = 22;
        end

         22 :
        begin                                                                   // tally
          //$display("AAAA %4d %4d tally", steps, ip);
            ip = 23;
        end

         23 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 24;
        end

         24 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 25;
              heapClock = ~ heapClock;
        end

         25 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[545] = heapOut;                                                     // Data retrieved from heap memory
              ip = 26;
              heapClock = ~ heapClock;
        end

         26 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[6] = localMem[545];
              ip = 27;
        end

         27 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[6] != 0 ? 79 : 28;
        end

         28 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 29;
              heapClock = ~ heapClock;
        end

         29 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[7] = heapOut;
              ip = 30;
        end

         30 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[546] = 1;
              ip = 31;
        end

         31 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[546];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 32;
              heapClock = ~ heapClock;
        end

         32 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[547] = 0;
              ip = 33;
        end

         33 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[547];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 34;
              heapClock = ~ heapClock;
        end

         34 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 35;
              heapClock = ~ heapClock;
        end

         35 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[8] = heapOut;
              ip = 36;
        end

         36 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[548] = localMem[8];
              ip = 37;
        end

         37 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[548];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 38;
              heapClock = ~ heapClock;
        end

         38 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 39;
              heapClock = ~ heapClock;
        end

         39 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[9] = heapOut;
              ip = 40;
        end

         40 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[549] = localMem[9];
              ip = 41;
        end

         41 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[549];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 42;
              heapClock = ~ heapClock;
        end

         42 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[550] = 0;
              ip = 43;
        end

         43 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[550];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 44;
              heapClock = ~ heapClock;
        end

         44 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[551] = localMem[0];
              ip = 45;
        end

         45 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[551];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 46;
              heapClock = ~ heapClock;
        end

         46 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 47;
              heapClock = ~ heapClock;
        end

         47 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[552] = heapOut;                                                     // Data retrieved from heap memory
              ip = 48;
              heapClock = ~ heapClock;
        end

         48 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[553] = localMem[552] + 1;
              ip = 49;
        end

         49 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[553];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 50;
              heapClock = ~ heapClock;
        end

         50 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 51;
              heapClock = ~ heapClock;
        end

         51 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[554] = heapOut;                                                     // Data retrieved from heap memory
              ip = 52;
              heapClock = ~ heapClock;
        end

         52 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[555] = localMem[554];
              ip = 53;
        end

         53 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[7];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[555];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 54;
              heapClock = ~ heapClock;
        end

         54 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[7];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 55;
              heapClock = ~ heapClock;
        end

         55 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[556] = heapOut;                                                     // Data retrieved from heap memory
              ip = 56;
              heapClock = ~ heapClock;
        end

         56 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[10] = localMem[556];
              ip = 57;
        end

         57 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[557] = localMem[3];
              ip = 58;
        end

         58 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[10];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[557];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 59;
              heapClock = ~ heapClock;
        end

         59 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[7];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 60;
              heapClock = ~ heapClock;
        end

         60 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[558] = heapOut;                                                     // Data retrieved from heap memory
              ip = 61;
              heapClock = ~ heapClock;
        end

         61 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[11] = localMem[558];
              ip = 62;
        end

         62 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[559] = localMem[5];
              ip = 63;
        end

         63 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[11];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[559];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 64;
              heapClock = ~ heapClock;
        end

         64 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 65;
              heapClock = ~ heapClock;
        end

         65 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[560] = heapOut;                                                     // Data retrieved from heap memory
              ip = 66;
              heapClock = ~ heapClock;
        end

         66 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[561] = localMem[560] + 1;
              ip = 67;
        end

         67 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[561];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 68;
              heapClock = ~ heapClock;
        end

         68 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[562] = localMem[7];
              ip = 69;
        end

         69 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[562];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 70;
              heapClock = ~ heapClock;
        end

         70 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[7];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 71;
              heapClock = ~ heapClock;
        end

         71 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[563] = heapOut;                                                     // Data retrieved from heap memory
              ip = 72;
              heapClock = ~ heapClock;
        end

         72 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[12] = localMem[563];
              ip = 73;
        end

         73 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[12];
              ip = 74;
              heapClock = ~ heapClock;
        end

         74 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[7];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 75;
              heapClock = ~ heapClock;
        end

         75 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[564] = heapOut;                                                     // Data retrieved from heap memory
              ip = 76;
              heapClock = ~ heapClock;
        end

         76 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[13] = localMem[564];
              ip = 77;
        end

         77 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[13];
              ip = 78;
              heapClock = ~ heapClock;
        end

         78 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2164;
        end

         79 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 80;
        end

         80 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 81;
              heapClock = ~ heapClock;
        end

         81 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[565] = heapOut;                                                     // Data retrieved from heap memory
              ip = 82;
              heapClock = ~ heapClock;
        end

         82 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[14] = localMem[565];
              ip = 83;
        end

         83 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 84;
              heapClock = ~ heapClock;
        end

         84 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[566] = heapOut;                                                     // Data retrieved from heap memory
              ip = 85;
              heapClock = ~ heapClock;
        end

         85 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[15] = localMem[566];
              ip = 86;
        end

         86 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[14] >= localMem[15] ? 156 : 87;
        end

         87 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 88;
              heapClock = ~ heapClock;
        end

         88 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[567] = heapOut;                                                     // Data retrieved from heap memory
              ip = 89;
              heapClock = ~ heapClock;
        end

         89 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[16] = localMem[567];
              ip = 90;
        end

         90 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[16] != 0 ? 155 : 91;
        end

         91 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 92;
              heapClock = ~ heapClock;
        end

         92 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[568] = heapOut;                                                     // Data retrieved from heap memory
              ip = 93;
              heapClock = ~ heapClock;
        end

         93 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[17] = !localMem[568];
              ip = 94;
        end

         94 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[17] == 0 ? 154 : 95;
        end

         95 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 96;
              heapClock = ~ heapClock;
        end

         96 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[569] = heapOut;                                                     // Data retrieved from heap memory
              ip = 97;
              heapClock = ~ heapClock;
        end

         97 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[18] = localMem[569];
              ip = 98;
        end

         98 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[3];
              heapAction = `Index;
              heapArray  = localMem[18];
              ip = 99;
              heapClock = ~ heapClock;
        end

         99 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[19] = heapOut;
              ip = 100;
        end

        100 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[19] == 0 ? 108 : 101;
        end

        101 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   101");
        end

        102 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   102");
        end

        103 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   103");
        end

        104 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   104");
        end

        105 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   105");
        end

        106 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   106");
        end

        107 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   107");
        end

        108 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 109;
        end

        109 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[14];
              heapArray  = localMem[18];
              ip = 110;
              heapClock = ~ heapClock;
        end

        110 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 111;
              heapClock = ~ heapClock;
        end

        111 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[572] = heapOut;                                                     // Data retrieved from heap memory
              ip = 112;
              heapClock = ~ heapClock;
        end

        112 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[21] = localMem[572];
              ip = 113;
        end

        113 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = localMem[14];
              heapArray  = localMem[21];
              ip = 114;
              heapClock = ~ heapClock;
        end

        114 :
        begin                                                                   // arrayCountGreater
          //$display("AAAA %4d %4d arrayCountGreater", steps, ip);
              heapIn     = localMem[3];
              heapAction = `Greater;
              heapArray  = localMem[18];
              ip = 115;
              heapClock = ~ heapClock;
        end

        115 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[22] = heapOut;
              ip = 116;
        end

        116 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[22] != 0 ? 134 : 117;
        end

        117 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 118;
              heapClock = ~ heapClock;
        end

        118 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[573] = heapOut;                                                     // Data retrieved from heap memory
              ip = 119;
              heapClock = ~ heapClock;
        end

        119 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[23] = localMem[573];
              ip = 120;
        end

        120 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[574] = localMem[3];
              ip = 121;
        end

        121 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[23];                                                // Array to write to
              heapIndex   = localMem[14];                                                // Index of element to write to
              heapIn      = localMem[574];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 122;
              heapClock = ~ heapClock;
        end

        122 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 123;
              heapClock = ~ heapClock;
        end

        123 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[575] = heapOut;                                                     // Data retrieved from heap memory
              ip = 124;
              heapClock = ~ heapClock;
        end

        124 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[24] = localMem[575];
              ip = 125;
        end

        125 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[576] = localMem[5];
              ip = 126;
        end

        126 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[24];                                                // Array to write to
              heapIndex   = localMem[14];                                                // Index of element to write to
              heapIn      = localMem[576];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 127;
              heapClock = ~ heapClock;
        end

        127 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[577] = localMem[14] + 1;
              ip = 128;
        end

        128 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[6];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[577];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 129;
              heapClock = ~ heapClock;
        end

        129 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 130;
              heapClock = ~ heapClock;
        end

        130 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[578] = heapOut;                                                     // Data retrieved from heap memory
              ip = 131;
              heapClock = ~ heapClock;
        end

        131 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[579] = localMem[578] + 1;
              ip = 132;
        end

        132 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[579];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 133;
              heapClock = ~ heapClock;
        end

        133 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2164;
        end

        134 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 135;
        end

        135 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
              heapIn     = localMem[3];
              heapAction = `Less;
              heapArray  = localMem[18];
              ip = 136;
              heapClock = ~ heapClock;
        end

        136 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[25] = heapOut;
              ip = 137;
        end

        137 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 138;
              heapClock = ~ heapClock;
        end

        138 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[580] = heapOut;                                                     // Data retrieved from heap memory
              ip = 139;
              heapClock = ~ heapClock;
        end

        139 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[26] = localMem[580];
              ip = 140;
        end

        140 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[3];
              heapArray  = localMem[26];
              heapIndex  = localMem[25];
              ip = 141;
              heapClock = ~ heapClock;
        end

        141 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 142;
              heapClock = ~ heapClock;
        end

        142 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[581] = heapOut;                                                     // Data retrieved from heap memory
              ip = 143;
              heapClock = ~ heapClock;
        end

        143 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[27] = localMem[581];
              ip = 144;
        end

        144 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[5];
              heapArray  = localMem[27];
              heapIndex  = localMem[25];
              ip = 145;
              heapClock = ~ heapClock;
        end

        145 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[6];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 146;
              heapClock = ~ heapClock;
        end

        146 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[582] = heapOut;                                                     // Data retrieved from heap memory
              ip = 147;
              heapClock = ~ heapClock;
        end

        147 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[583] = localMem[582] + 1;
              ip = 148;
        end

        148 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[6];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[583];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 149;
              heapClock = ~ heapClock;
        end

        149 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 150;
              heapClock = ~ heapClock;
        end

        150 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[584] = heapOut;                                                     // Data retrieved from heap memory
              ip = 151;
              heapClock = ~ heapClock;
        end

        151 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[585] = localMem[584] + 1;
              ip = 152;
        end

        152 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[585];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 153;
              heapClock = ~ heapClock;
        end

        153 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2164;
        end

        154 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 155;
        end

        155 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 156;
        end

        156 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 157;
        end

        157 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 158;
              heapClock = ~ heapClock;
        end

        158 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[586] = heapOut;                                                     // Data retrieved from heap memory
              ip = 159;
              heapClock = ~ heapClock;
        end

        159 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[28] = localMem[586];
              ip = 160;
        end

        160 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 161;
        end

        161 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 162;
              heapClock = ~ heapClock;
        end

        162 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[587] = heapOut;                                                     // Data retrieved from heap memory
              ip = 163;
              heapClock = ~ heapClock;
        end

        163 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[30] = localMem[587];
              ip = 164;
        end

        164 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[30] <  3 ? 624 : 165;
        end

        165 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 166;
              heapClock = ~ heapClock;
        end

        166 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[588] = heapOut;                                                     // Data retrieved from heap memory
              ip = 167;
              heapClock = ~ heapClock;
        end

        167 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[31] = localMem[588];
              ip = 168;
        end

        168 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 169;
              heapClock = ~ heapClock;
        end

        169 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[589] = heapOut;                                                     // Data retrieved from heap memory
              ip = 170;
              heapClock = ~ heapClock;
        end

        170 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[32] = localMem[589];
              ip = 171;
        end

        171 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[32] == 0 ? 375 : 172;
        end

        172 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   172");
        end

        173 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   173");
        end

        174 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   174");
        end

        175 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   175");
        end

        176 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   176");
        end

        177 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   177");
        end

        178 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   178");
        end

        179 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   179");
        end

        180 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   180");
        end

        181 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   181");
        end

        182 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   182");
        end

        183 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   183");
        end

        184 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   184");
        end

        185 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   185");
        end

        186 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   186");
        end

        187 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   187");
        end

        188 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   188");
        end

        189 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   189");
        end

        190 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   190");
        end

        191 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   191");
        end

        192 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   192");
        end

        193 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   193");
        end

        194 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   194");
        end

        195 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   195");
        end

        196 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   196");
        end

        197 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   197");
        end

        198 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   198");
        end

        199 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   199");
        end

        200 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   200");
        end

        201 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   201");
        end

        202 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   202");
        end

        203 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   203");
        end

        204 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   204");
        end

        205 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   205");
        end

        206 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   206");
        end

        207 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   207");
        end

        208 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   208");
        end

        209 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   209");
        end

        210 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   210");
        end

        211 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   211");
        end

        212 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   212");
        end

        213 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   213");
        end

        214 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   214");
        end

        215 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   215");
        end

        216 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   216");
        end

        217 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   217");
        end

        218 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   218");
        end

        219 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   219");
        end

        220 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   220");
        end

        221 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   221");
        end

        222 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   222");
        end

        223 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   223");
        end

        224 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   224");
        end

        225 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   225");
        end

        226 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   226");
        end

        227 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   227");
        end

        228 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   228");
        end

        229 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   229");
        end

        230 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   230");
        end

        231 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   231");
        end

        232 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   232");
        end

        233 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   233");
        end

        234 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   234");
        end

        235 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   235");
        end

        236 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   236");
        end

        237 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   237");
        end

        238 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   238");
        end

        239 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   239");
        end

        240 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   240");
        end

        241 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed   241");
        end

        242 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   242");
        end

        243 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   243");
        end

        244 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   244");
        end

        245 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   245");
        end

        246 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   246");
        end

        247 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   247");
        end

        248 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   248");
        end

        249 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   249");
        end

        250 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   250");
        end

        251 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   251");
        end

        252 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   252");
        end

        253 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   253");
        end

        254 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   254");
        end

        255 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   255");
        end

        256 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   256");
        end

        257 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   257");
        end

        258 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   258");
        end

        259 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   259");
        end

        260 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   260");
        end

        261 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   261");
        end

        262 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   262");
        end

        263 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   263");
        end

        264 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   264");
        end

        265 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   265");
        end

        266 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   266");
        end

        267 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   267");
        end

        268 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   268");
        end

        269 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   269");
        end

        270 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   270");
        end

        271 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   271");
        end

        272 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   272");
        end

        273 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   273");
        end

        274 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   274");
        end

        275 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   275");
        end

        276 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   276");
        end

        277 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   277");
        end

        278 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   278");
        end

        279 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   279");
        end

        280 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   280");
        end

        281 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   281");
        end

        282 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   282");
        end

        283 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   283");
        end

        284 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   284");
        end

        285 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   285");
        end

        286 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   286");
        end

        287 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   287");
        end

        288 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   288");
        end

        289 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   289");
        end

        290 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   290");
        end

        291 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   291");
        end

        292 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   292");
        end

        293 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   293");
        end

        294 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   294");
        end

        295 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   295");
        end

        296 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   296");
        end

        297 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   297");
        end

        298 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   298");
        end

        299 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   299");
        end

        300 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   300");
        end

        301 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   301");
        end

        302 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   302");
        end

        303 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   303");
        end

        304 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   304");
        end

        305 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   305");
        end

        306 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   306");
        end

        307 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   307");
        end

        308 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   308");
        end

        309 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   309");
        end

        310 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   310");
        end

        311 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   311");
        end

        312 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   312");
        end

        313 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   313");
        end

        314 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   314");
        end

        315 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   315");
        end

        316 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   316");
        end

        317 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   317");
        end

        318 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   318");
        end

        319 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   319");
        end

        320 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   320");
        end

        321 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   321");
        end

        322 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   322");
        end

        323 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   323");
        end

        324 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   324");
        end

        325 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   325");
        end

        326 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   326");
        end

        327 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   327");
        end

        328 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   328");
        end

        329 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   329");
        end

        330 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   330");
        end

        331 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   331");
        end

        332 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   332");
        end

        333 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   333");
        end

        334 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   334");
        end

        335 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   335");
        end

        336 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   336");
        end

        337 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   337");
        end

        338 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   338");
        end

        339 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   339");
        end

        340 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   340");
        end

        341 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   341");
        end

        342 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   342");
        end

        343 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   343");
        end

        344 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   344");
        end

        345 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   345");
        end

        346 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   346");
        end

        347 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   347");
        end

        348 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   348");
        end

        349 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   349");
        end

        350 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   350");
        end

        351 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   351");
        end

        352 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   352");
        end

        353 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   353");
        end

        354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   354");
        end

        355 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   355");
        end

        356 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   356");
        end

        357 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   357");
        end

        358 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   358");
        end

        359 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   359");
        end

        360 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   360");
        end

        361 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   361");
        end

        362 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   362");
        end

        363 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   363");
        end

        364 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   364");
        end

        365 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   365");
        end

        366 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   366");
        end

        367 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   367");
        end

        368 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   368");
        end

        369 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   369");
        end

        370 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   370");
        end

        371 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   371");
        end

        372 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   372");
        end

        373 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   373");
        end

        374 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   374");
        end

        375 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 376;
        end

        376 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 377;
              heapClock = ~ heapClock;
        end

        377 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[80] = heapOut;
              ip = 378;
        end

        378 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[647] = 1;
              ip = 379;
        end

        379 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[647];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 380;
              heapClock = ~ heapClock;
        end

        380 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[648] = 0;
              ip = 381;
        end

        381 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[648];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 382;
              heapClock = ~ heapClock;
        end

        382 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 383;
              heapClock = ~ heapClock;
        end

        383 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[81] = heapOut;
              ip = 384;
        end

        384 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[649] = localMem[81];
              ip = 385;
        end

        385 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[649];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 386;
              heapClock = ~ heapClock;
        end

        386 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 387;
              heapClock = ~ heapClock;
        end

        387 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[82] = heapOut;
              ip = 388;
        end

        388 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[650] = localMem[82];
              ip = 389;
        end

        389 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[650];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 390;
              heapClock = ~ heapClock;
        end

        390 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[651] = 0;
              ip = 391;
        end

        391 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[651];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 392;
              heapClock = ~ heapClock;
        end

        392 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[652] = localMem[31];
              ip = 393;
        end

        393 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[652];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 394;
              heapClock = ~ heapClock;
        end

        394 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 395;
              heapClock = ~ heapClock;
        end

        395 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[653] = heapOut;                                                     // Data retrieved from heap memory
              ip = 396;
              heapClock = ~ heapClock;
        end

        396 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[654] = localMem[653] + 1;
              ip = 397;
        end

        397 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[31];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[654];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 398;
              heapClock = ~ heapClock;
        end

        398 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 399;
              heapClock = ~ heapClock;
        end

        399 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[655] = heapOut;                                                     // Data retrieved from heap memory
              ip = 400;
              heapClock = ~ heapClock;
        end

        400 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[656] = localMem[655];
              ip = 401;
        end

        401 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[656];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 402;
              heapClock = ~ heapClock;
        end

        402 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 403;
              heapClock = ~ heapClock;
        end

        403 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[83] = heapOut;
              ip = 404;
        end

        404 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[657] = 1;
              ip = 405;
        end

        405 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[657];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 406;
              heapClock = ~ heapClock;
        end

        406 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[658] = 0;
              ip = 407;
        end

        407 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[658];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 408;
              heapClock = ~ heapClock;
        end

        408 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 409;
              heapClock = ~ heapClock;
        end

        409 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[84] = heapOut;
              ip = 410;
        end

        410 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[659] = localMem[84];
              ip = 411;
        end

        411 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[659];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 412;
              heapClock = ~ heapClock;
        end

        412 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 413;
              heapClock = ~ heapClock;
        end

        413 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[85] = heapOut;
              ip = 414;
        end

        414 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[660] = localMem[85];
              ip = 415;
        end

        415 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[660];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 416;
              heapClock = ~ heapClock;
        end

        416 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[661] = 0;
              ip = 417;
        end

        417 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[661];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 418;
              heapClock = ~ heapClock;
        end

        418 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[662] = localMem[31];
              ip = 419;
        end

        419 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[662];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 420;
              heapClock = ~ heapClock;
        end

        420 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 421;
              heapClock = ~ heapClock;
        end

        421 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[663] = heapOut;                                                     // Data retrieved from heap memory
              ip = 422;
              heapClock = ~ heapClock;
        end

        422 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[664] = localMem[663] + 1;
              ip = 423;
        end

        423 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[31];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[664];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 424;
              heapClock = ~ heapClock;
        end

        424 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[31];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 425;
              heapClock = ~ heapClock;
        end

        425 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[665] = heapOut;                                                     // Data retrieved from heap memory
              ip = 426;
              heapClock = ~ heapClock;
        end

        426 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[666] = localMem[665];
              ip = 427;
        end

        427 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[666];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 428;
              heapClock = ~ heapClock;
        end

        428 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 429;
              heapClock = ~ heapClock;
        end

        429 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[667] = heapOut;                                                     // Data retrieved from heap memory
              ip = 430;
              heapClock = ~ heapClock;
        end

        430 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[86] = !localMem[667];
              ip = 431;
        end

        431 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[86] != 0 ? 531 : 432;
        end

        432 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 433;
              heapClock = ~ heapClock;
        end

        433 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[87] = heapOut;
              ip = 434;
        end

        434 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[668] = localMem[87];
              ip = 435;
        end

        435 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[668];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 436;
              heapClock = ~ heapClock;
        end

        436 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 437;
              heapClock = ~ heapClock;
        end

        437 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[88] = heapOut;
              ip = 438;
        end

        438 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[669] = localMem[88];
              ip = 439;
        end

        439 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[669];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 440;
              heapClock = ~ heapClock;
        end

        440 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 441;
              heapClock = ~ heapClock;
        end

        441 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[670] = heapOut;                                                     // Data retrieved from heap memory
              ip = 442;
              heapClock = ~ heapClock;
        end

        442 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[89] = localMem[670];
              ip = 443;
        end

        443 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[80];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 444;
              heapClock = ~ heapClock;
        end

        444 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[671] = heapOut;                                                     // Data retrieved from heap memory
              ip = 445;
              heapClock = ~ heapClock;
        end

        445 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[90] = localMem[671];
              ip = 446;
        end

        446 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[89];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 447;
              heapClock = ~ heapClock;
        end

        447 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[90];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 448;
              heapClock = ~ heapClock;
        end

        448 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 449;
              heapClock = ~ heapClock;
        end

        449 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[672] = heapOut;                                                     // Data retrieved from heap memory
              ip = 450;
              heapClock = ~ heapClock;
        end

        450 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[91] = localMem[672];
              ip = 451;
        end

        451 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[80];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 452;
              heapClock = ~ heapClock;
        end

        452 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[673] = heapOut;                                                     // Data retrieved from heap memory
              ip = 453;
              heapClock = ~ heapClock;
        end

        453 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[92] = localMem[673];
              ip = 454;
        end

        454 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[91];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 455;
              heapClock = ~ heapClock;
        end

        455 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[92];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 456;
              heapClock = ~ heapClock;
        end

        456 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 457;
              heapClock = ~ heapClock;
        end

        457 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[674] = heapOut;                                                     // Data retrieved from heap memory
              ip = 458;
              heapClock = ~ heapClock;
        end

        458 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[93] = localMem[674];
              ip = 459;
        end

        459 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[80];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 460;
              heapClock = ~ heapClock;
        end

        460 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[675] = heapOut;                                                     // Data retrieved from heap memory
              ip = 461;
              heapClock = ~ heapClock;
        end

        461 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[94] = localMem[675];
              ip = 462;
        end

        462 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[95] = 1 + 1;
              ip = 463;
        end

        463 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[93];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 464;
              heapClock = ~ heapClock;
        end

        464 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[94];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[95];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 465;
              heapClock = ~ heapClock;
        end

        465 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 466;
              heapClock = ~ heapClock;
        end

        466 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[676] = heapOut;                                                     // Data retrieved from heap memory
              ip = 467;
              heapClock = ~ heapClock;
        end

        467 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[96] = localMem[676];
              ip = 468;
        end

        468 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[83];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 469;
              heapClock = ~ heapClock;
        end

        469 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[677] = heapOut;                                                     // Data retrieved from heap memory
              ip = 470;
              heapClock = ~ heapClock;
        end

        470 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[97] = localMem[677];
              ip = 471;
        end

        471 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[96];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 472;
              heapClock = ~ heapClock;
        end

        472 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[97];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 473;
              heapClock = ~ heapClock;
        end

        473 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 474;
              heapClock = ~ heapClock;
        end

        474 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[678] = heapOut;                                                     // Data retrieved from heap memory
              ip = 475;
              heapClock = ~ heapClock;
        end

        475 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[98] = localMem[678];
              ip = 476;
        end

        476 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[83];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 477;
              heapClock = ~ heapClock;
        end

        477 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[679] = heapOut;                                                     // Data retrieved from heap memory
              ip = 478;
              heapClock = ~ heapClock;
        end

        478 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[99] = localMem[679];
              ip = 479;
        end

        479 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[98];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 480;
              heapClock = ~ heapClock;
        end

        480 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[99];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 481;
              heapClock = ~ heapClock;
        end

        481 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 482;
              heapClock = ~ heapClock;
        end

        482 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[680] = heapOut;                                                     // Data retrieved from heap memory
              ip = 483;
              heapClock = ~ heapClock;
        end

        483 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[100] = localMem[680];
              ip = 484;
        end

        484 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[83];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 485;
              heapClock = ~ heapClock;
        end

        485 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[681] = heapOut;                                                     // Data retrieved from heap memory
              ip = 486;
              heapClock = ~ heapClock;
        end

        486 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[101] = localMem[681];
              ip = 487;
        end

        487 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[102] = 1 + 1;
              ip = 488;
        end

        488 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[100];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 489;
              heapClock = ~ heapClock;
        end

        489 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[101];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[102];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 490;
              heapClock = ~ heapClock;
        end

        490 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[80];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 491;
              heapClock = ~ heapClock;
        end

        491 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[682] = heapOut;                                                     // Data retrieved from heap memory
              ip = 492;
              heapClock = ~ heapClock;
        end

        492 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[103] = localMem[682];
              ip = 493;
        end

        493 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[104] = localMem[103] + 1;
              ip = 494;
        end

        494 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[80];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 495;
              heapClock = ~ heapClock;
        end

        495 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[683] = heapOut;                                                     // Data retrieved from heap memory
              ip = 496;
              heapClock = ~ heapClock;
        end

        496 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[105] = localMem[683];
              ip = 497;
        end

        497 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 498;
        end

        498 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[106] = 0;
              ip = 499;
        end

        499 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 500;
        end

        500 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[106] >= localMem[104] ? 509 : 501;
        end

        501 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[105];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[106];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 502;
              heapClock = ~ heapClock;
        end

        502 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[684] = heapOut;                                                     // Data retrieved from heap memory
              ip = 503;
              heapClock = ~ heapClock;
        end

        503 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[107] = localMem[684];
              ip = 504;
        end

        504 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[685] = localMem[80];
              ip = 505;
        end

        505 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[107];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[685];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 506;
              heapClock = ~ heapClock;
        end

        506 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 507;
        end

        507 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[106] = localMem[106] + 1;
              ip = 508;
        end

        508 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 499;
        end

        509 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 510;
        end

        510 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[83];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 511;
              heapClock = ~ heapClock;
        end

        511 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[686] = heapOut;                                                     // Data retrieved from heap memory
              ip = 512;
              heapClock = ~ heapClock;
        end

        512 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[108] = localMem[686];
              ip = 513;
        end

        513 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[109] = localMem[108] + 1;
              ip = 514;
        end

        514 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[83];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 515;
              heapClock = ~ heapClock;
        end

        515 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[687] = heapOut;                                                     // Data retrieved from heap memory
              ip = 516;
              heapClock = ~ heapClock;
        end

        516 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[110] = localMem[687];
              ip = 517;
        end

        517 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 518;
        end

        518 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[111] = 0;
              ip = 519;
        end

        519 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 520;
        end

        520 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[111] >= localMem[109] ? 529 : 521;
        end

        521 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[110];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[111];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 522;
              heapClock = ~ heapClock;
        end

        522 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[688] = heapOut;                                                     // Data retrieved from heap memory
              ip = 523;
              heapClock = ~ heapClock;
        end

        523 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[112] = localMem[688];
              ip = 524;
        end

        524 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[689] = localMem[83];
              ip = 525;
        end

        525 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[112];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[689];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 526;
              heapClock = ~ heapClock;
        end

        526 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 527;
        end

        527 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[111] = localMem[111] + 1;
              ip = 528;
        end

        528 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 519;
        end

        529 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 530;
        end

        530 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 568;
        end

        531 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 532;
        end

        532 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 533;
              heapClock = ~ heapClock;
        end

        533 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[113] = heapOut;
              ip = 534;
        end

        534 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[690] = localMem[113];
              ip = 535;
        end

        535 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[28];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[690];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 536;
              heapClock = ~ heapClock;
        end

        536 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 537;
              heapClock = ~ heapClock;
        end

        537 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[691] = heapOut;                                                     // Data retrieved from heap memory
              ip = 538;
              heapClock = ~ heapClock;
        end

        538 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[114] = localMem[691];
              ip = 539;
        end

        539 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[80];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 540;
              heapClock = ~ heapClock;
        end

        540 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[692] = heapOut;                                                     // Data retrieved from heap memory
              ip = 541;
              heapClock = ~ heapClock;
        end

        541 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[115] = localMem[692];
              ip = 542;
        end

        542 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[114];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 543;
              heapClock = ~ heapClock;
        end

        543 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[115];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 544;
              heapClock = ~ heapClock;
        end

        544 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 545;
              heapClock = ~ heapClock;
        end

        545 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[693] = heapOut;                                                     // Data retrieved from heap memory
              ip = 546;
              heapClock = ~ heapClock;
        end

        546 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[116] = localMem[693];
              ip = 547;
        end

        547 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[80];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 548;
              heapClock = ~ heapClock;
        end

        548 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[694] = heapOut;                                                     // Data retrieved from heap memory
              ip = 549;
              heapClock = ~ heapClock;
        end

        549 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[117] = localMem[694];
              ip = 550;
        end

        550 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[116];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 551;
              heapClock = ~ heapClock;
        end

        551 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[117];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 552;
              heapClock = ~ heapClock;
        end

        552 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 553;
              heapClock = ~ heapClock;
        end

        553 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[695] = heapOut;                                                     // Data retrieved from heap memory
              ip = 554;
              heapClock = ~ heapClock;
        end

        554 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[118] = localMem[695];
              ip = 555;
        end

        555 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[83];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 556;
              heapClock = ~ heapClock;
        end

        556 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[696] = heapOut;                                                     // Data retrieved from heap memory
              ip = 557;
              heapClock = ~ heapClock;
        end

        557 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[119] = localMem[696];
              ip = 558;
        end

        558 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[118];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 559;
              heapClock = ~ heapClock;
        end

        559 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[119];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 560;
              heapClock = ~ heapClock;
        end

        560 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 561;
              heapClock = ~ heapClock;
        end

        561 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[697] = heapOut;                                                     // Data retrieved from heap memory
              ip = 562;
              heapClock = ~ heapClock;
        end

        562 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[120] = localMem[697];
              ip = 563;
        end

        563 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[83];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 564;
              heapClock = ~ heapClock;
        end

        564 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[698] = heapOut;                                                     // Data retrieved from heap memory
              ip = 565;
              heapClock = ~ heapClock;
        end

        565 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[121] = localMem[698];
              ip = 566;
        end

        566 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[120];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 567;
              heapClock = ~ heapClock;
        end

        567 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[121];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 568;
              heapClock = ~ heapClock;
        end

        568 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 569;
        end

        569 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[699] = localMem[28];
              ip = 570;
        end

        570 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[80];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[699];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 571;
              heapClock = ~ heapClock;
        end

        571 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[700] = localMem[28];
              ip = 572;
        end

        572 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[83];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[700];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 573;
              heapClock = ~ heapClock;
        end

        573 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 574;
              heapClock = ~ heapClock;
        end

        574 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[701] = heapOut;                                                     // Data retrieved from heap memory
              ip = 575;
              heapClock = ~ heapClock;
        end

        575 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[122] = localMem[701];
              ip = 576;
        end

        576 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[122];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 577;
              heapClock = ~ heapClock;
        end

        577 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[702] = heapOut;                                                     // Data retrieved from heap memory
              ip = 578;
              heapClock = ~ heapClock;
        end

        578 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[123] = localMem[702];
              ip = 579;
        end

        579 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 580;
              heapClock = ~ heapClock;
        end

        580 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[703] = heapOut;                                                     // Data retrieved from heap memory
              ip = 581;
              heapClock = ~ heapClock;
        end

        581 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[124] = localMem[703];
              ip = 582;
        end

        582 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[124];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 583;
              heapClock = ~ heapClock;
        end

        583 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[704] = heapOut;                                                     // Data retrieved from heap memory
              ip = 584;
              heapClock = ~ heapClock;
        end

        584 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[125] = localMem[704];
              ip = 585;
        end

        585 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 586;
              heapClock = ~ heapClock;
        end

        586 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[705] = heapOut;                                                     // Data retrieved from heap memory
              ip = 587;
              heapClock = ~ heapClock;
        end

        587 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[126] = localMem[705];
              ip = 588;
        end

        588 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[706] = localMem[123];
              ip = 589;
        end

        589 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[126];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[706];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 590;
              heapClock = ~ heapClock;
        end

        590 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 591;
              heapClock = ~ heapClock;
        end

        591 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[707] = heapOut;                                                     // Data retrieved from heap memory
              ip = 592;
              heapClock = ~ heapClock;
        end

        592 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[127] = localMem[707];
              ip = 593;
        end

        593 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[708] = localMem[125];
              ip = 594;
        end

        594 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[127];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[708];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 595;
              heapClock = ~ heapClock;
        end

        595 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 596;
              heapClock = ~ heapClock;
        end

        596 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[709] = heapOut;                                                     // Data retrieved from heap memory
              ip = 597;
              heapClock = ~ heapClock;
        end

        597 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[128] = localMem[709];
              ip = 598;
        end

        598 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[710] = localMem[80];
              ip = 599;
        end

        599 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[128];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[710];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 600;
              heapClock = ~ heapClock;
        end

        600 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 601;
              heapClock = ~ heapClock;
        end

        601 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[711] = heapOut;                                                     // Data retrieved from heap memory
              ip = 602;
              heapClock = ~ heapClock;
        end

        602 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[129] = localMem[711];
              ip = 603;
        end

        603 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[712] = localMem[83];
              ip = 604;
        end

        604 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[129];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[712];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 605;
              heapClock = ~ heapClock;
        end

        605 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[713] = 1;
              ip = 606;
        end

        606 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[28];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[713];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 607;
              heapClock = ~ heapClock;
        end

        607 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 608;
              heapClock = ~ heapClock;
        end

        608 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[714] = heapOut;                                                     // Data retrieved from heap memory
              ip = 609;
              heapClock = ~ heapClock;
        end

        609 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[130] = localMem[714];
              ip = 610;
        end

        610 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[130];
              ip = 611;
              heapClock = ~ heapClock;
        end

        611 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 612;
              heapClock = ~ heapClock;
        end

        612 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[715] = heapOut;                                                     // Data retrieved from heap memory
              ip = 613;
              heapClock = ~ heapClock;
        end

        613 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[131] = localMem[715];
              ip = 614;
        end

        614 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[131];
              ip = 615;
              heapClock = ~ heapClock;
        end

        615 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 616;
              heapClock = ~ heapClock;
        end

        616 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[716] = heapOut;                                                     // Data retrieved from heap memory
              ip = 617;
              heapClock = ~ heapClock;
        end

        617 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[132] = localMem[716];
              ip = 618;
        end

        618 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 2;
              heapArray  = localMem[132];
              ip = 619;
              heapClock = ~ heapClock;
        end

        619 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 621;
        end

        620 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   620");
        end

        621 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 622;
        end

        622 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[29] = 1;
              ip = 623;
        end

        623 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 626;
        end

        624 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 625;
        end

        625 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[29] = 0;
              ip = 626;
        end

        626 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 627;
        end

        627 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 628;
        end

        628 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 629;
        end

        629 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[133] = 0;
              ip = 630;
        end

        630 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 631;
        end

        631 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[133] >= 99 ? 1640 : 632;
        end

        632 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 633;
              heapClock = ~ heapClock;
        end

        633 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[717] = heapOut;                                                     // Data retrieved from heap memory
              ip = 634;
              heapClock = ~ heapClock;
        end

        634 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[134] = localMem[717];
              ip = 635;
        end

        635 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[135] = localMem[134] - 1;
              ip = 636;
        end

        636 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 637;
              heapClock = ~ heapClock;
        end

        637 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[718] = heapOut;                                                     // Data retrieved from heap memory
              ip = 638;
              heapClock = ~ heapClock;
        end

        638 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[136] = localMem[718];
              ip = 639;
        end

        639 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[136];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[135];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 640;
              heapClock = ~ heapClock;
        end

        640 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[719] = heapOut;                                                     // Data retrieved from heap memory
              ip = 641;
              heapClock = ~ heapClock;
        end

        641 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[137] = localMem[719];
              ip = 642;
        end

        642 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[3] <= localMem[137] ? 1132 : 643;
        end

        643 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 644;
              heapClock = ~ heapClock;
        end

        644 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[720] = heapOut;                                                     // Data retrieved from heap memory
              ip = 645;
              heapClock = ~ heapClock;
        end

        645 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[138] = !localMem[720];
              ip = 646;
        end

        646 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[138] == 0 ? 654 : 647;
        end

        647 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[721] = localMem[28];
              ip = 648;
        end

        648 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[721];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 649;
              heapClock = ~ heapClock;
        end

        649 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[722] = 2;
              ip = 650;
        end

        650 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[722];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 651;
              heapClock = ~ heapClock;
        end

        651 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[723] = localMem[134] - 1;
              ip = 652;
        end

        652 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[723];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 653;
              heapClock = ~ heapClock;
        end

        653 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1644;
        end

        654 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 655;
        end

        655 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 656;
              heapClock = ~ heapClock;
        end

        656 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[724] = heapOut;                                                     // Data retrieved from heap memory
              ip = 657;
              heapClock = ~ heapClock;
        end

        657 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[139] = localMem[724];
              ip = 658;
        end

        658 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[139];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[134];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 659;
              heapClock = ~ heapClock;
        end

        659 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[725] = heapOut;                                                     // Data retrieved from heap memory
              ip = 660;
              heapClock = ~ heapClock;
        end

        660 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[140] = localMem[725];
              ip = 661;
        end

        661 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 662;
        end

        662 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 663;
              heapClock = ~ heapClock;
        end

        663 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[726] = heapOut;                                                     // Data retrieved from heap memory
              ip = 664;
              heapClock = ~ heapClock;
        end

        664 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[142] = localMem[726];
              ip = 665;
        end

        665 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[142] <  3 ? 1125 : 666;
        end

        666 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 667;
              heapClock = ~ heapClock;
        end

        667 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[727] = heapOut;                                                     // Data retrieved from heap memory
              ip = 668;
              heapClock = ~ heapClock;
        end

        668 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[143] = localMem[727];
              ip = 669;
        end

        669 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 670;
              heapClock = ~ heapClock;
        end

        670 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[728] = heapOut;                                                     // Data retrieved from heap memory
              ip = 671;
              heapClock = ~ heapClock;
        end

        671 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[144] = localMem[728];
              ip = 672;
        end

        672 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[144] == 0 ? 876 : 673;
        end

        673 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 674;
              heapClock = ~ heapClock;
        end

        674 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[145] = heapOut;
              ip = 675;
        end

        675 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[729] = 1;
              ip = 676;
        end

        676 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[729];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 677;
              heapClock = ~ heapClock;
        end

        677 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[730] = 0;
              ip = 678;
        end

        678 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[730];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 679;
              heapClock = ~ heapClock;
        end

        679 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 680;
              heapClock = ~ heapClock;
        end

        680 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[146] = heapOut;
              ip = 681;
        end

        681 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[731] = localMem[146];
              ip = 682;
        end

        682 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[731];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 683;
              heapClock = ~ heapClock;
        end

        683 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 684;
              heapClock = ~ heapClock;
        end

        684 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[147] = heapOut;
              ip = 685;
        end

        685 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[732] = localMem[147];
              ip = 686;
        end

        686 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[732];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 687;
              heapClock = ~ heapClock;
        end

        687 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[733] = 0;
              ip = 688;
        end

        688 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[733];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 689;
              heapClock = ~ heapClock;
        end

        689 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[734] = localMem[143];
              ip = 690;
        end

        690 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[734];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 691;
              heapClock = ~ heapClock;
        end

        691 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[143];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 692;
              heapClock = ~ heapClock;
        end

        692 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[735] = heapOut;                                                     // Data retrieved from heap memory
              ip = 693;
              heapClock = ~ heapClock;
        end

        693 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[736] = localMem[735] + 1;
              ip = 694;
        end

        694 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[143];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[736];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 695;
              heapClock = ~ heapClock;
        end

        695 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[143];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 696;
              heapClock = ~ heapClock;
        end

        696 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[737] = heapOut;                                                     // Data retrieved from heap memory
              ip = 697;
              heapClock = ~ heapClock;
        end

        697 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[738] = localMem[737];
              ip = 698;
        end

        698 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[738];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 699;
              heapClock = ~ heapClock;
        end

        699 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 700;
              heapClock = ~ heapClock;
        end

        700 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[739] = heapOut;                                                     // Data retrieved from heap memory
              ip = 701;
              heapClock = ~ heapClock;
        end

        701 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[148] = !localMem[739];
              ip = 702;
        end

        702 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[148] != 0 ? 757 : 703;
        end

        703 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 704;
              heapClock = ~ heapClock;
        end

        704 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[149] = heapOut;
              ip = 705;
        end

        705 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[740] = localMem[149];
              ip = 706;
        end

        706 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[740];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 707;
              heapClock = ~ heapClock;
        end

        707 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 708;
              heapClock = ~ heapClock;
        end

        708 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[741] = heapOut;                                                     // Data retrieved from heap memory
              ip = 709;
              heapClock = ~ heapClock;
        end

        709 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[150] = localMem[741];
              ip = 710;
        end

        710 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[145];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 711;
              heapClock = ~ heapClock;
        end

        711 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[742] = heapOut;                                                     // Data retrieved from heap memory
              ip = 712;
              heapClock = ~ heapClock;
        end

        712 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[151] = localMem[742];
              ip = 713;
        end

        713 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[150];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 714;
              heapClock = ~ heapClock;
        end

        714 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[151];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 715;
              heapClock = ~ heapClock;
        end

        715 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 716;
              heapClock = ~ heapClock;
        end

        716 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[743] = heapOut;                                                     // Data retrieved from heap memory
              ip = 717;
              heapClock = ~ heapClock;
        end

        717 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[152] = localMem[743];
              ip = 718;
        end

        718 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[145];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 719;
              heapClock = ~ heapClock;
        end

        719 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[744] = heapOut;                                                     // Data retrieved from heap memory
              ip = 720;
              heapClock = ~ heapClock;
        end

        720 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[153] = localMem[744];
              ip = 721;
        end

        721 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[152];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 722;
              heapClock = ~ heapClock;
        end

        722 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[153];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 723;
              heapClock = ~ heapClock;
        end

        723 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 724;
              heapClock = ~ heapClock;
        end

        724 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[745] = heapOut;                                                     // Data retrieved from heap memory
              ip = 725;
              heapClock = ~ heapClock;
        end

        725 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[154] = localMem[745];
              ip = 726;
        end

        726 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[145];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 727;
              heapClock = ~ heapClock;
        end

        727 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[746] = heapOut;                                                     // Data retrieved from heap memory
              ip = 728;
              heapClock = ~ heapClock;
        end

        728 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[155] = localMem[746];
              ip = 729;
        end

        729 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[156] = 1 + 1;
              ip = 730;
        end

        730 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[154];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 731;
              heapClock = ~ heapClock;
        end

        731 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[155];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[156];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 732;
              heapClock = ~ heapClock;
        end

        732 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[145];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 733;
              heapClock = ~ heapClock;
        end

        733 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[747] = heapOut;                                                     // Data retrieved from heap memory
              ip = 734;
              heapClock = ~ heapClock;
        end

        734 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[157] = localMem[747];
              ip = 735;
        end

        735 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[158] = localMem[157] + 1;
              ip = 736;
        end

        736 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[145];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 737;
              heapClock = ~ heapClock;
        end

        737 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[748] = heapOut;                                                     // Data retrieved from heap memory
              ip = 738;
              heapClock = ~ heapClock;
        end

        738 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[159] = localMem[748];
              ip = 739;
        end

        739 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 740;
        end

        740 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[160] = 0;
              ip = 741;
        end

        741 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 742;
        end

        742 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[160] >= localMem[158] ? 751 : 743;
        end

        743 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[159];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[160];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 744;
              heapClock = ~ heapClock;
        end

        744 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[749] = heapOut;                                                     // Data retrieved from heap memory
              ip = 745;
              heapClock = ~ heapClock;
        end

        745 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[161] = localMem[749];
              ip = 746;
        end

        746 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[750] = localMem[145];
              ip = 747;
        end

        747 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[161];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[750];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 748;
              heapClock = ~ heapClock;
        end

        748 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 749;
        end

        749 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[160] = localMem[160] + 1;
              ip = 750;
        end

        750 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 741;
        end

        751 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 752;
        end

        752 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 753;
              heapClock = ~ heapClock;
        end

        753 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[751] = heapOut;                                                     // Data retrieved from heap memory
              ip = 754;
              heapClock = ~ heapClock;
        end

        754 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[162] = localMem[751];
              ip = 755;
        end

        755 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 2;
              heapArray  = localMem[162];
              ip = 756;
              heapClock = ~ heapClock;
        end

        756 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 774;
        end

        757 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   757");
        end

        758 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   758");
        end

        759 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   759");
        end

        760 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   760");
        end

        761 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   761");
        end

        762 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   762");
        end

        763 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   763");
        end

        764 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   764");
        end

        765 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   765");
        end

        766 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   766");
        end

        767 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   767");
        end

        768 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   768");
        end

        769 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   769");
        end

        770 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   770");
        end

        771 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   771");
        end

        772 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   772");
        end

        773 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   773");
        end

        774 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 775;
        end

        775 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[756] = 1;
              ip = 776;
        end

        776 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[140];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[756];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 777;
              heapClock = ~ heapClock;
        end

        777 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[757] = localMem[144];
              ip = 778;
        end

        778 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[145];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[757];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 779;
              heapClock = ~ heapClock;
        end

        779 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 780;
              heapClock = ~ heapClock;
        end

        780 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[758] = heapOut;                                                     // Data retrieved from heap memory
              ip = 781;
              heapClock = ~ heapClock;
        end

        781 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[167] = localMem[758];
              ip = 782;
        end

        782 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 783;
              heapClock = ~ heapClock;
        end

        783 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[759] = heapOut;                                                     // Data retrieved from heap memory
              ip = 784;
              heapClock = ~ heapClock;
        end

        784 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[168] = localMem[759];
              ip = 785;
        end

        785 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[168];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[167];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 786;
              heapClock = ~ heapClock;
        end

        786 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[760] = heapOut;                                                     // Data retrieved from heap memory
              ip = 787;
              heapClock = ~ heapClock;
        end

        787 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[169] = localMem[760];
              ip = 788;
        end

        788 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[169] != localMem[140] ? 829 : 789;
        end

        789 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 790;
              heapClock = ~ heapClock;
        end

        790 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[761] = heapOut;                                                     // Data retrieved from heap memory
              ip = 791;
              heapClock = ~ heapClock;
        end

        791 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[170] = localMem[761];
              ip = 792;
        end

        792 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[170];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 793;
              heapClock = ~ heapClock;
        end

        793 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[762] = heapOut;                                                     // Data retrieved from heap memory
              ip = 794;
              heapClock = ~ heapClock;
        end

        794 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[171] = localMem[762];
              ip = 795;
        end

        795 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 796;
              heapClock = ~ heapClock;
        end

        796 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[763] = heapOut;                                                     // Data retrieved from heap memory
              ip = 797;
              heapClock = ~ heapClock;
        end

        797 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[172] = localMem[763];
              ip = 798;
        end

        798 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[764] = localMem[171];
              ip = 799;
        end

        799 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[172];                                                // Array to write to
              heapIndex   = localMem[167];                                                // Index of element to write to
              heapIn      = localMem[764];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 800;
              heapClock = ~ heapClock;
        end

        800 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 801;
              heapClock = ~ heapClock;
        end

        801 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[765] = heapOut;                                                     // Data retrieved from heap memory
              ip = 802;
              heapClock = ~ heapClock;
        end

        802 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[173] = localMem[765];
              ip = 803;
        end

        803 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[173];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 804;
              heapClock = ~ heapClock;
        end

        804 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[766] = heapOut;                                                     // Data retrieved from heap memory
              ip = 805;
              heapClock = ~ heapClock;
        end

        805 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[174] = localMem[766];
              ip = 806;
        end

        806 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 807;
              heapClock = ~ heapClock;
        end

        807 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[767] = heapOut;                                                     // Data retrieved from heap memory
              ip = 808;
              heapClock = ~ heapClock;
        end

        808 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[175] = localMem[767];
              ip = 809;
        end

        809 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[768] = localMem[174];
              ip = 810;
        end

        810 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[175];                                                // Array to write to
              heapIndex   = localMem[167];                                                // Index of element to write to
              heapIn      = localMem[768];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 811;
              heapClock = ~ heapClock;
        end

        811 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 812;
              heapClock = ~ heapClock;
        end

        812 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[769] = heapOut;                                                     // Data retrieved from heap memory
              ip = 813;
              heapClock = ~ heapClock;
        end

        813 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[176] = localMem[769];
              ip = 814;
        end

        814 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[176];
              ip = 815;
              heapClock = ~ heapClock;
        end

        815 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[140];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 816;
              heapClock = ~ heapClock;
        end

        816 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[770] = heapOut;                                                     // Data retrieved from heap memory
              ip = 817;
              heapClock = ~ heapClock;
        end

        817 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[177] = localMem[770];
              ip = 818;
        end

        818 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[177];
              ip = 819;
              heapClock = ~ heapClock;
        end

        819 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[178] = localMem[167] + 1;
              ip = 820;
        end

        820 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[771] = localMem[178];
              ip = 821;
        end

        821 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[144];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[771];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 822;
              heapClock = ~ heapClock;
        end

        822 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[144];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 823;
              heapClock = ~ heapClock;
        end

        823 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[772] = heapOut;                                                     // Data retrieved from heap memory
              ip = 824;
              heapClock = ~ heapClock;
        end

        824 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[179] = localMem[772];
              ip = 825;
        end

        825 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[773] = localMem[145];
              ip = 826;
        end

        826 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[179];                                                // Array to write to
              heapIndex   = localMem[178];                                                // Index of element to write to
              heapIn      = localMem[773];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 827;
              heapClock = ~ heapClock;
        end

        827 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1122;
        end

        828 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   828");
        end

        829 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   829");
        end

        830 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
          // $display("Should not be executed   830");
        end

        831 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   831");
        end

        832 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   832");
        end

        833 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   833");
        end

        834 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
          // $display("Should not be executed   834");
        end

        835 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   835");
        end

        836 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed   836");
        end

        837 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   837");
        end

        838 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   838");
        end

        839 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   839");
        end

        840 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   840");
        end

        841 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   841");
        end

        842 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   842");
        end

        843 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   843");
        end

        844 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   844");
        end

        845 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   845");
        end

        846 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   846");
        end

        847 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   847");
        end

        848 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   848");
        end

        849 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   849");
        end

        850 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   850");
        end

        851 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   851");
        end

        852 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   852");
        end

        853 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   853");
        end

        854 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   854");
        end

        855 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   855");
        end

        856 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed   856");
        end

        857 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   857");
        end

        858 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   858");
        end

        859 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   859");
        end

        860 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   860");
        end

        861 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   861");
        end

        862 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   862");
        end

        863 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   863");
        end

        864 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   864");
        end

        865 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   865");
        end

        866 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   866");
        end

        867 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   867");
        end

        868 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   868");
        end

        869 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
          // $display("Should not be executed   869");
        end

        870 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   870");
        end

        871 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   871");
        end

        872 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   872");
        end

        873 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   873");
        end

        874 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed   874");
        end

        875 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   875");
        end

        876 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   876");
        end

        877 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   877");
        end

        878 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   878");
        end

        879 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   879");
        end

        880 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   880");
        end

        881 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   881");
        end

        882 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   882");
        end

        883 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   883");
        end

        884 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   884");
        end

        885 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   885");
        end

        886 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   886");
        end

        887 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   887");
        end

        888 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   888");
        end

        889 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   889");
        end

        890 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   890");
        end

        891 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   891");
        end

        892 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   892");
        end

        893 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   893");
        end

        894 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   894");
        end

        895 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   895");
        end

        896 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   896");
        end

        897 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   897");
        end

        898 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   898");
        end

        899 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   899");
        end

        900 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   900");
        end

        901 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   901");
        end

        902 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   902");
        end

        903 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   903");
        end

        904 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   904");
        end

        905 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   905");
        end

        906 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   906");
        end

        907 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   907");
        end

        908 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   908");
        end

        909 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   909");
        end

        910 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   910");
        end

        911 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   911");
        end

        912 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   912");
        end

        913 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   913");
        end

        914 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   914");
        end

        915 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   915");
        end

        916 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   916");
        end

        917 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   917");
        end

        918 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   918");
        end

        919 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   919");
        end

        920 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   920");
        end

        921 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   921");
        end

        922 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   922");
        end

        923 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   923");
        end

        924 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   924");
        end

        925 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   925");
        end

        926 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   926");
        end

        927 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   927");
        end

        928 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   928");
        end

        929 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   929");
        end

        930 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   930");
        end

        931 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed   931");
        end

        932 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed   932");
        end

        933 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   933");
        end

        934 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   934");
        end

        935 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   935");
        end

        936 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   936");
        end

        937 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed   937");
        end

        938 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed   938");
        end

        939 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   939");
        end

        940 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed   940");
        end

        941 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   941");
        end

        942 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   942");
        end

        943 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   943");
        end

        944 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   944");
        end

        945 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   945");
        end

        946 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   946");
        end

        947 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   947");
        end

        948 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   948");
        end

        949 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   949");
        end

        950 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   950");
        end

        951 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   951");
        end

        952 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   952");
        end

        953 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   953");
        end

        954 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   954");
        end

        955 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   955");
        end

        956 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   956");
        end

        957 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   957");
        end

        958 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   958");
        end

        959 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   959");
        end

        960 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   960");
        end

        961 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   961");
        end

        962 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   962");
        end

        963 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   963");
        end

        964 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   964");
        end

        965 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   965");
        end

        966 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   966");
        end

        967 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   967");
        end

        968 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   968");
        end

        969 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   969");
        end

        970 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   970");
        end

        971 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   971");
        end

        972 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   972");
        end

        973 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   973");
        end

        974 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   974");
        end

        975 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   975");
        end

        976 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   976");
        end

        977 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   977");
        end

        978 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   978");
        end

        979 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   979");
        end

        980 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   980");
        end

        981 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   981");
        end

        982 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   982");
        end

        983 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   983");
        end

        984 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   984");
        end

        985 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   985");
        end

        986 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   986");
        end

        987 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   987");
        end

        988 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   988");
        end

        989 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed   989");
        end

        990 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed   990");
        end

        991 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   991");
        end

        992 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   992");
        end

        993 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   993");
        end

        994 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed   994");
        end

        995 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed   995");
        end

        996 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed   996");
        end

        997 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   997");
        end

        998 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed   998");
        end

        999 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed   999");
        end

       1000 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1000");
        end

       1001 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1001");
        end

       1002 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1002");
        end

       1003 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1003");
        end

       1004 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1004");
        end

       1005 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1005");
        end

       1006 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1006");
        end

       1007 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1007");
        end

       1008 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1008");
        end

       1009 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1009");
        end

       1010 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1010");
        end

       1011 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1011");
        end

       1012 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1012");
        end

       1013 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1013");
        end

       1014 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1014");
        end

       1015 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1015");
        end

       1016 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1016");
        end

       1017 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1017");
        end

       1018 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1018");
        end

       1019 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1019");
        end

       1020 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1020");
        end

       1021 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1021");
        end

       1022 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1022");
        end

       1023 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1023");
        end

       1024 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1024");
        end

       1025 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1025");
        end

       1026 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1026");
        end

       1027 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1027");
        end

       1028 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1028");
        end

       1029 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1029");
        end

       1030 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1030");
        end

       1031 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1031");
        end

       1032 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1032");
        end

       1033 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1033");
        end

       1034 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1034");
        end

       1035 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1035");
        end

       1036 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1036");
        end

       1037 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1037");
        end

       1038 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1038");
        end

       1039 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1039");
        end

       1040 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1040");
        end

       1041 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1041");
        end

       1042 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1042");
        end

       1043 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1043");
        end

       1044 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1044");
        end

       1045 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1045");
        end

       1046 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1046");
        end

       1047 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1047");
        end

       1048 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1048");
        end

       1049 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1049");
        end

       1050 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1050");
        end

       1051 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1051");
        end

       1052 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1052");
        end

       1053 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1053");
        end

       1054 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1054");
        end

       1055 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1055");
        end

       1056 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1056");
        end

       1057 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1057");
        end

       1058 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1058");
        end

       1059 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1059");
        end

       1060 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1060");
        end

       1061 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1061");
        end

       1062 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1062");
        end

       1063 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1063");
        end

       1064 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1064");
        end

       1065 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1065");
        end

       1066 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1066");
        end

       1067 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1067");
        end

       1068 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1068");
        end

       1069 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1069");
        end

       1070 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1070");
        end

       1071 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1071");
        end

       1072 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1072");
        end

       1073 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1073");
        end

       1074 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1074");
        end

       1075 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1075");
        end

       1076 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1076");
        end

       1077 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1077");
        end

       1078 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1078");
        end

       1079 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1079");
        end

       1080 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1080");
        end

       1081 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1081");
        end

       1082 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1082");
        end

       1083 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1083");
        end

       1084 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1084");
        end

       1085 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1085");
        end

       1086 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1086");
        end

       1087 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1087");
        end

       1088 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1088");
        end

       1089 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1089");
        end

       1090 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1090");
        end

       1091 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1091");
        end

       1092 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1092");
        end

       1093 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1093");
        end

       1094 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1094");
        end

       1095 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1095");
        end

       1096 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1096");
        end

       1097 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1097");
        end

       1098 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1098");
        end

       1099 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1099");
        end

       1100 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1100");
        end

       1101 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1101");
        end

       1102 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1102");
        end

       1103 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1103");
        end

       1104 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1104");
        end

       1105 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1105");
        end

       1106 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1106");
        end

       1107 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1107");
        end

       1108 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1108");
        end

       1109 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1109");
        end

       1110 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1110");
        end

       1111 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1111");
        end

       1112 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1112");
        end

       1113 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1113");
        end

       1114 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1114");
        end

       1115 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1115");
        end

       1116 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1116");
        end

       1117 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1117");
        end

       1118 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1118");
        end

       1119 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1119");
        end

       1120 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1120");
        end

       1121 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1121");
        end

       1122 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1123;
        end

       1123 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[141] = 1;
              ip = 1124;
        end

       1124 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1127;
        end

       1125 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1126;
        end

       1126 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[141] = 0;
              ip = 1127;
        end

       1127 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1128;
        end

       1128 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[141] != 0 ? 1130 : 1129;
        end

       1129 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[28] = localMem[140];
              ip = 1130;
        end

       1130 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1131;
        end

       1131 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1637;
        end

       1132 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1133;
        end

       1133 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1134;
              heapClock = ~ heapClock;
        end

       1134 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[856] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1135;
              heapClock = ~ heapClock;
        end

       1135 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[245] = localMem[856];
              ip = 1136;
        end

       1136 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[3];
              heapAction = `Index;
              heapArray  = localMem[245];
              ip = 1137;
              heapClock = ~ heapClock;
        end

       1137 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[246] = heapOut;
              ip = 1138;
        end

       1138 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[246] == 0 ? 1146 : 1139;
        end

       1139 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1139");
        end

       1140 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1140");
        end

       1141 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1141");
        end

       1142 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1142");
        end

       1143 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
          // $display("Should not be executed  1143");
        end

       1144 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1144");
        end

       1145 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1145");
        end

       1146 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1147;
        end

       1147 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
              heapIn     = localMem[3];
              heapAction = `Less;
              heapArray  = localMem[245];
              ip = 1148;
              heapClock = ~ heapClock;
        end

       1148 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[247] = heapOut;
              ip = 1149;
        end

       1149 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1150;
              heapClock = ~ heapClock;
        end

       1150 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[860] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1151;
              heapClock = ~ heapClock;
        end

       1151 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[248] = !localMem[860];
              ip = 1152;
        end

       1152 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[248] == 0 ? 1160 : 1153;
        end

       1153 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[861] = localMem[28];
              ip = 1154;
        end

       1154 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[861];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1155;
              heapClock = ~ heapClock;
        end

       1155 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[862] = 0;
              ip = 1156;
        end

       1156 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[862];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1157;
              heapClock = ~ heapClock;
        end

       1157 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[863] = localMem[247];
              ip = 1158;
        end

       1158 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[863];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1159;
              heapClock = ~ heapClock;
        end

       1159 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1644;
        end

       1160 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1161;
        end

       1161 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[28];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1162;
              heapClock = ~ heapClock;
        end

       1162 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[864] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1163;
              heapClock = ~ heapClock;
        end

       1163 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[249] = localMem[864];
              ip = 1164;
        end

       1164 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[249];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[247];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1165;
              heapClock = ~ heapClock;
        end

       1165 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[865] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1166;
              heapClock = ~ heapClock;
        end

       1166 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[250] = localMem[865];
              ip = 1167;
        end

       1167 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1168;
        end

       1168 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1169;
              heapClock = ~ heapClock;
        end

       1169 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[866] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1170;
              heapClock = ~ heapClock;
        end

       1170 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[252] = localMem[866];
              ip = 1171;
        end

       1171 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[252] <  3 ? 1631 : 1172;
        end

       1172 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1173;
              heapClock = ~ heapClock;
        end

       1173 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[867] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1174;
              heapClock = ~ heapClock;
        end

       1174 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[253] = localMem[867];
              ip = 1175;
        end

       1175 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1176;
              heapClock = ~ heapClock;
        end

       1176 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[868] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1177;
              heapClock = ~ heapClock;
        end

       1177 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[254] = localMem[868];
              ip = 1178;
        end

       1178 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[254] == 0 ? 1382 : 1179;
        end

       1179 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1180;
              heapClock = ~ heapClock;
        end

       1180 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[255] = heapOut;
              ip = 1181;
        end

       1181 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[869] = 1;
              ip = 1182;
        end

       1182 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[869];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1183;
              heapClock = ~ heapClock;
        end

       1183 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[870] = 0;
              ip = 1184;
        end

       1184 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[870];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1185;
              heapClock = ~ heapClock;
        end

       1185 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1186;
              heapClock = ~ heapClock;
        end

       1186 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[256] = heapOut;
              ip = 1187;
        end

       1187 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[871] = localMem[256];
              ip = 1188;
        end

       1188 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[871];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1189;
              heapClock = ~ heapClock;
        end

       1189 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1190;
              heapClock = ~ heapClock;
        end

       1190 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[257] = heapOut;
              ip = 1191;
        end

       1191 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[872] = localMem[257];
              ip = 1192;
        end

       1192 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[872];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1193;
              heapClock = ~ heapClock;
        end

       1193 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[873] = 0;
              ip = 1194;
        end

       1194 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[873];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1195;
              heapClock = ~ heapClock;
        end

       1195 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[874] = localMem[253];
              ip = 1196;
        end

       1196 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[874];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1197;
              heapClock = ~ heapClock;
        end

       1197 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[253];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1198;
              heapClock = ~ heapClock;
        end

       1198 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[875] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1199;
              heapClock = ~ heapClock;
        end

       1199 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[876] = localMem[875] + 1;
              ip = 1200;
        end

       1200 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[253];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[876];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1201;
              heapClock = ~ heapClock;
        end

       1201 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[253];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1202;
              heapClock = ~ heapClock;
        end

       1202 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[877] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1203;
              heapClock = ~ heapClock;
        end

       1203 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[878] = localMem[877];
              ip = 1204;
        end

       1204 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[878];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1205;
              heapClock = ~ heapClock;
        end

       1205 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1206;
              heapClock = ~ heapClock;
        end

       1206 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[879] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1207;
              heapClock = ~ heapClock;
        end

       1207 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[258] = !localMem[879];
              ip = 1208;
        end

       1208 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[258] != 0 ? 1263 : 1209;
        end

       1209 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1210;
              heapClock = ~ heapClock;
        end

       1210 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[259] = heapOut;
              ip = 1211;
        end

       1211 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[880] = localMem[259];
              ip = 1212;
        end

       1212 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[880];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1213;
              heapClock = ~ heapClock;
        end

       1213 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1214;
              heapClock = ~ heapClock;
        end

       1214 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[881] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1215;
              heapClock = ~ heapClock;
        end

       1215 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[260] = localMem[881];
              ip = 1216;
        end

       1216 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[255];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1217;
              heapClock = ~ heapClock;
        end

       1217 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[882] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1218;
              heapClock = ~ heapClock;
        end

       1218 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[261] = localMem[882];
              ip = 1219;
        end

       1219 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[260];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1220;
              heapClock = ~ heapClock;
        end

       1220 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[261];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1221;
              heapClock = ~ heapClock;
        end

       1221 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1222;
              heapClock = ~ heapClock;
        end

       1222 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[883] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1223;
              heapClock = ~ heapClock;
        end

       1223 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[262] = localMem[883];
              ip = 1224;
        end

       1224 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[255];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1225;
              heapClock = ~ heapClock;
        end

       1225 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[884] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1226;
              heapClock = ~ heapClock;
        end

       1226 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[263] = localMem[884];
              ip = 1227;
        end

       1227 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[262];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1228;
              heapClock = ~ heapClock;
        end

       1228 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[263];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1229;
              heapClock = ~ heapClock;
        end

       1229 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1230;
              heapClock = ~ heapClock;
        end

       1230 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[885] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1231;
              heapClock = ~ heapClock;
        end

       1231 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[264] = localMem[885];
              ip = 1232;
        end

       1232 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[255];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1233;
              heapClock = ~ heapClock;
        end

       1233 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[886] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1234;
              heapClock = ~ heapClock;
        end

       1234 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[265] = localMem[886];
              ip = 1235;
        end

       1235 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[266] = 1 + 1;
              ip = 1236;
        end

       1236 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[264];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1237;
              heapClock = ~ heapClock;
        end

       1237 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[265];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = localMem[266];                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1238;
              heapClock = ~ heapClock;
        end

       1238 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[255];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1239;
              heapClock = ~ heapClock;
        end

       1239 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[887] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1240;
              heapClock = ~ heapClock;
        end

       1240 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[267] = localMem[887];
              ip = 1241;
        end

       1241 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[268] = localMem[267] + 1;
              ip = 1242;
        end

       1242 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[255];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1243;
              heapClock = ~ heapClock;
        end

       1243 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[888] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1244;
              heapClock = ~ heapClock;
        end

       1244 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[269] = localMem[888];
              ip = 1245;
        end

       1245 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1246;
        end

       1246 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[270] = 0;
              ip = 1247;
        end

       1247 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1248;
        end

       1248 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[270] >= localMem[268] ? 1257 : 1249;
        end

       1249 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[269];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[270];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1250;
              heapClock = ~ heapClock;
        end

       1250 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[889] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1251;
              heapClock = ~ heapClock;
        end

       1251 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[271] = localMem[889];
              ip = 1252;
        end

       1252 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[890] = localMem[255];
              ip = 1253;
        end

       1253 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[271];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[890];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1254;
              heapClock = ~ heapClock;
        end

       1254 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1255;
        end

       1255 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[270] = localMem[270] + 1;
              ip = 1256;
        end

       1256 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1247;
        end

       1257 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1258;
        end

       1258 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1259;
              heapClock = ~ heapClock;
        end

       1259 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[891] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1260;
              heapClock = ~ heapClock;
        end

       1260 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[272] = localMem[891];
              ip = 1261;
        end

       1261 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 2;
              heapArray  = localMem[272];
              ip = 1262;
              heapClock = ~ heapClock;
        end

       1262 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1280;
        end

       1263 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1263");
        end

       1264 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1264");
        end

       1265 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1265");
        end

       1266 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1266");
        end

       1267 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1267");
        end

       1268 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1268");
        end

       1269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1269");
        end

       1270 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1270");
        end

       1271 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1271");
        end

       1272 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1272");
        end

       1273 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1273");
        end

       1274 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1274");
        end

       1275 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1275");
        end

       1276 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1276");
        end

       1277 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1277");
        end

       1278 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1278");
        end

       1279 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1279");
        end

       1280 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1281;
        end

       1281 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[896] = 1;
              ip = 1282;
        end

       1282 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[250];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[896];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1283;
              heapClock = ~ heapClock;
        end

       1283 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[897] = localMem[254];
              ip = 1284;
        end

       1284 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[255];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[897];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1285;
              heapClock = ~ heapClock;
        end

       1285 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[254];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1286;
              heapClock = ~ heapClock;
        end

       1286 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[898] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1287;
              heapClock = ~ heapClock;
        end

       1287 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[277] = localMem[898];
              ip = 1288;
        end

       1288 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[254];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1289;
              heapClock = ~ heapClock;
        end

       1289 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[899] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1290;
              heapClock = ~ heapClock;
        end

       1290 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[278] = localMem[899];
              ip = 1291;
        end

       1291 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[278];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[277];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1292;
              heapClock = ~ heapClock;
        end

       1292 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[900] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1293;
              heapClock = ~ heapClock;
        end

       1293 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[279] = localMem[900];
              ip = 1294;
        end

       1294 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[279] != localMem[250] ? 1335 : 1295;
        end

       1295 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1295");
        end

       1296 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1296");
        end

       1297 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1297");
        end

       1298 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1298");
        end

       1299 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1299");
        end

       1300 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1300");
        end

       1301 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1301");
        end

       1302 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1302");
        end

       1303 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1303");
        end

       1304 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1304");
        end

       1305 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1305");
        end

       1306 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1306");
        end

       1307 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1307");
        end

       1308 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1308");
        end

       1309 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1309");
        end

       1310 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1310");
        end

       1311 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1311");
        end

       1312 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1312");
        end

       1313 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1313");
        end

       1314 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1314");
        end

       1315 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1315");
        end

       1316 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1316");
        end

       1317 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1317");
        end

       1318 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1318");
        end

       1319 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1319");
        end

       1320 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1320");
        end

       1321 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1321");
        end

       1322 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1322");
        end

       1323 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1323");
        end

       1324 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1324");
        end

       1325 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1325");
        end

       1326 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1326");
        end

       1327 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1327");
        end

       1328 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1328");
        end

       1329 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1329");
        end

       1330 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1330");
        end

       1331 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1331");
        end

       1332 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1332");
        end

       1333 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1333");
        end

       1334 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1334");
        end

       1335 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1336;
        end

       1336 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
            ip = 1337;
        end

       1337 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[254];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1338;
              heapClock = ~ heapClock;
        end

       1338 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[914] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1339;
              heapClock = ~ heapClock;
        end

       1339 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[290] = localMem[914];
              ip = 1340;
        end

       1340 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[250];
              heapAction = `Index;
              heapArray  = localMem[290];
              ip = 1341;
              heapClock = ~ heapClock;
        end

       1341 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[291] = heapOut;
              ip = 1342;
        end

       1342 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[291] = localMem[291] - 1;
              ip = 1343;
        end

       1343 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1344;
              heapClock = ~ heapClock;
        end

       1344 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[915] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1345;
              heapClock = ~ heapClock;
        end

       1345 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[292] = localMem[915];
              ip = 1346;
        end

       1346 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[292];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1347;
              heapClock = ~ heapClock;
        end

       1347 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[916] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1348;
              heapClock = ~ heapClock;
        end

       1348 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[293] = localMem[916];
              ip = 1349;
        end

       1349 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1350;
              heapClock = ~ heapClock;
        end

       1350 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[917] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1351;
              heapClock = ~ heapClock;
        end

       1351 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[294] = localMem[917];
              ip = 1352;
        end

       1352 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[294];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1353;
              heapClock = ~ heapClock;
        end

       1353 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[918] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1354;
              heapClock = ~ heapClock;
        end

       1354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[295] = localMem[918];
              ip = 1355;
        end

       1355 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1356;
              heapClock = ~ heapClock;
        end

       1356 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[919] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1357;
              heapClock = ~ heapClock;
        end

       1357 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[296] = localMem[919];
              ip = 1358;
        end

       1358 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[296];
              ip = 1359;
              heapClock = ~ heapClock;
        end

       1359 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[250];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1360;
              heapClock = ~ heapClock;
        end

       1360 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[920] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1361;
              heapClock = ~ heapClock;
        end

       1361 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[297] = localMem[920];
              ip = 1362;
        end

       1362 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[297];
              ip = 1363;
              heapClock = ~ heapClock;
        end

       1363 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[254];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1364;
              heapClock = ~ heapClock;
        end

       1364 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[921] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1365;
              heapClock = ~ heapClock;
        end

       1365 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[298] = localMem[921];
              ip = 1366;
        end

       1366 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[293];
              heapArray  = localMem[298];
              heapIndex  = localMem[291];
              ip = 1367;
              heapClock = ~ heapClock;
        end

       1367 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[254];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1368;
              heapClock = ~ heapClock;
        end

       1368 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[922] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1369;
              heapClock = ~ heapClock;
        end

       1369 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[299] = localMem[922];
              ip = 1370;
        end

       1370 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[295];
              heapArray  = localMem[299];
              heapIndex  = localMem[291];
              ip = 1371;
              heapClock = ~ heapClock;
        end

       1371 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[254];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1372;
              heapClock = ~ heapClock;
        end

       1372 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[923] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1373;
              heapClock = ~ heapClock;
        end

       1373 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[300] = localMem[923];
              ip = 1374;
        end

       1374 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[301] = localMem[291] + 1;
              ip = 1375;
        end

       1375 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[255];
              heapArray  = localMem[300];
              heapIndex  = localMem[301];
              ip = 1376;
              heapClock = ~ heapClock;
        end

       1376 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[254];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1377;
              heapClock = ~ heapClock;
        end

       1377 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[924] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1378;
              heapClock = ~ heapClock;
        end

       1378 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[925] = localMem[924] + 1;
              ip = 1379;
        end

       1379 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[254];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[925];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1380;
              heapClock = ~ heapClock;
        end

       1380 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1628;
        end

       1381 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1381");
        end

       1382 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1382");
        end

       1383 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1383");
        end

       1384 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1384");
        end

       1385 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1385");
        end

       1386 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1386");
        end

       1387 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1387");
        end

       1388 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1388");
        end

       1389 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1389");
        end

       1390 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1390");
        end

       1391 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1391");
        end

       1392 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1392");
        end

       1393 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1393");
        end

       1394 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1394");
        end

       1395 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1395");
        end

       1396 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1396");
        end

       1397 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1397");
        end

       1398 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1398");
        end

       1399 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1399");
        end

       1400 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1400");
        end

       1401 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1401");
        end

       1402 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1402");
        end

       1403 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1403");
        end

       1404 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1404");
        end

       1405 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1405");
        end

       1406 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1406");
        end

       1407 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1407");
        end

       1408 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1408");
        end

       1409 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1409");
        end

       1410 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1410");
        end

       1411 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1411");
        end

       1412 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1412");
        end

       1413 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1413");
        end

       1414 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1414");
        end

       1415 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1415");
        end

       1416 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1416");
        end

       1417 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1417");
        end

       1418 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1418");
        end

       1419 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1419");
        end

       1420 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1420");
        end

       1421 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1421");
        end

       1422 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1422");
        end

       1423 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1423");
        end

       1424 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1424");
        end

       1425 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1425");
        end

       1426 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1426");
        end

       1427 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1427");
        end

       1428 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1428");
        end

       1429 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1429");
        end

       1430 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1430");
        end

       1431 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1431");
        end

       1432 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1432");
        end

       1433 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1433");
        end

       1434 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1434");
        end

       1435 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1435");
        end

       1436 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1436");
        end

       1437 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1437");
        end

       1438 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1438");
        end

       1439 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1439");
        end

       1440 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1440");
        end

       1441 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1441");
        end

       1442 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1442");
        end

       1443 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1443");
        end

       1444 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1444");
        end

       1445 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1445");
        end

       1446 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1446");
        end

       1447 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1447");
        end

       1448 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1448");
        end

       1449 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1449");
        end

       1450 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1450");
        end

       1451 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1451");
        end

       1452 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1452");
        end

       1453 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1453");
        end

       1454 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1454");
        end

       1455 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1455");
        end

       1456 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1456");
        end

       1457 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1457");
        end

       1458 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1458");
        end

       1459 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1459");
        end

       1460 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1460");
        end

       1461 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1461");
        end

       1462 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1462");
        end

       1463 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1463");
        end

       1464 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1464");
        end

       1465 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1465");
        end

       1466 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1466");
        end

       1467 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1467");
        end

       1468 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1468");
        end

       1469 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1469");
        end

       1470 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1470");
        end

       1471 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1471");
        end

       1472 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1472");
        end

       1473 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1473");
        end

       1474 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1474");
        end

       1475 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1475");
        end

       1476 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1476");
        end

       1477 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1477");
        end

       1478 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1478");
        end

       1479 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1479");
        end

       1480 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1480");
        end

       1481 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1481");
        end

       1482 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1482");
        end

       1483 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1483");
        end

       1484 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1484");
        end

       1485 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1485");
        end

       1486 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1486");
        end

       1487 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1487");
        end

       1488 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1488");
        end

       1489 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1489");
        end

       1490 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1490");
        end

       1491 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1491");
        end

       1492 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1492");
        end

       1493 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1493");
        end

       1494 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1494");
        end

       1495 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1495");
        end

       1496 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1496");
        end

       1497 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1497");
        end

       1498 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1498");
        end

       1499 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1499");
        end

       1500 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1500");
        end

       1501 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1501");
        end

       1502 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1502");
        end

       1503 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1503");
        end

       1504 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1504");
        end

       1505 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1505");
        end

       1506 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1506");
        end

       1507 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1507");
        end

       1508 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1508");
        end

       1509 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1509");
        end

       1510 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1510");
        end

       1511 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1511");
        end

       1512 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1512");
        end

       1513 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1513");
        end

       1514 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1514");
        end

       1515 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1515");
        end

       1516 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1516");
        end

       1517 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1517");
        end

       1518 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1518");
        end

       1519 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1519");
        end

       1520 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1520");
        end

       1521 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1521");
        end

       1522 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1522");
        end

       1523 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1523");
        end

       1524 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1524");
        end

       1525 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1525");
        end

       1526 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1526");
        end

       1527 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1527");
        end

       1528 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1528");
        end

       1529 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1529");
        end

       1530 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1530");
        end

       1531 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1531");
        end

       1532 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1532");
        end

       1533 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1533");
        end

       1534 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1534");
        end

       1535 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1535");
        end

       1536 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1536");
        end

       1537 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1537");
        end

       1538 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1538");
        end

       1539 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1539");
        end

       1540 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1540");
        end

       1541 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1541");
        end

       1542 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1542");
        end

       1543 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1543");
        end

       1544 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1544");
        end

       1545 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1545");
        end

       1546 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1546");
        end

       1547 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1547");
        end

       1548 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1548");
        end

       1549 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1549");
        end

       1550 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1550");
        end

       1551 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1551");
        end

       1552 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1552");
        end

       1553 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1553");
        end

       1554 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1554");
        end

       1555 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1555");
        end

       1556 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1556");
        end

       1557 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1557");
        end

       1558 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1558");
        end

       1559 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1559");
        end

       1560 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1560");
        end

       1561 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1561");
        end

       1562 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1562");
        end

       1563 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1563");
        end

       1564 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1564");
        end

       1565 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1565");
        end

       1566 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1566");
        end

       1567 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1567");
        end

       1568 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1568");
        end

       1569 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1569");
        end

       1570 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1570");
        end

       1571 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1571");
        end

       1572 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1572");
        end

       1573 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1573");
        end

       1574 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1574");
        end

       1575 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1575");
        end

       1576 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1576");
        end

       1577 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1577");
        end

       1578 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1578");
        end

       1579 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1579");
        end

       1580 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1580");
        end

       1581 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1581");
        end

       1582 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1582");
        end

       1583 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1583");
        end

       1584 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1584");
        end

       1585 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1585");
        end

       1586 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1586");
        end

       1587 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1587");
        end

       1588 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1588");
        end

       1589 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1589");
        end

       1590 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1590");
        end

       1591 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1591");
        end

       1592 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1592");
        end

       1593 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1593");
        end

       1594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1594");
        end

       1595 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1595");
        end

       1596 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1596");
        end

       1597 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1597");
        end

       1598 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1598");
        end

       1599 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1599");
        end

       1600 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1600");
        end

       1601 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1601");
        end

       1602 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1602");
        end

       1603 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1603");
        end

       1604 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1604");
        end

       1605 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1605");
        end

       1606 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1606");
        end

       1607 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1607");
        end

       1608 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1608");
        end

       1609 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1609");
        end

       1610 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1610");
        end

       1611 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1611");
        end

       1612 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1612");
        end

       1613 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1613");
        end

       1614 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1614");
        end

       1615 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1615");
        end

       1616 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1616");
        end

       1617 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1617");
        end

       1618 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1618");
        end

       1619 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1619");
        end

       1620 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1620");
        end

       1621 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1621");
        end

       1622 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1622");
        end

       1623 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1623");
        end

       1624 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1624");
        end

       1625 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1625");
        end

       1626 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1626");
        end

       1627 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1627");
        end

       1628 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1629;
        end

       1629 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[251] = 1;
              ip = 1630;
        end

       1630 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1633;
        end

       1631 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1632;
        end

       1632 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[251] = 0;
              ip = 1633;
        end

       1633 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1634;
        end

       1634 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[251] != 0 ? 1636 : 1635;
        end

       1635 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[28] = localMem[250];
              ip = 1636;
        end

       1636 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1637;
        end

       1637 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1638;
        end

       1638 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[133] = localMem[133] + 1;
              ip = 1639;
        end

       1639 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 630;
        end

       1640 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1640");
        end

       1641 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  1641");
        end

       1642 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1642");
        end

       1643 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1643");
        end

       1644 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1645;
        end

       1645 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[1];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1646;
              heapClock = ~ heapClock;
        end

       1646 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[996] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1647;
              heapClock = ~ heapClock;
        end

       1647 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[355] = localMem[996];
              ip = 1648;
        end

       1648 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[1];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1649;
              heapClock = ~ heapClock;
        end

       1649 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[997] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1650;
              heapClock = ~ heapClock;
        end

       1650 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[356] = localMem[997];
              ip = 1651;
        end

       1651 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[1];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1652;
              heapClock = ~ heapClock;
        end

       1652 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[998] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1653;
              heapClock = ~ heapClock;
        end

       1653 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[357] = localMem[998];
              ip = 1654;
        end

       1654 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[356] != 1 ? 1661 : 1655;
        end

       1655 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1655");
        end

       1656 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1656");
        end

       1657 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1657");
        end

       1658 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1658");
        end

       1659 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1659");
        end

       1660 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1660");
        end

       1661 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1662;
        end

       1662 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[356] != 2 ? 1677 : 1663;
        end

       1663 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[359] = localMem[357] + 1;
              ip = 1664;
        end

       1664 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1665;
              heapClock = ~ heapClock;
        end

       1665 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1001] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1666;
              heapClock = ~ heapClock;
        end

       1666 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[360] = localMem[1001];
              ip = 1667;
        end

       1667 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[3];
              heapArray  = localMem[360];
              heapIndex  = localMem[359];
              ip = 1668;
              heapClock = ~ heapClock;
        end

       1668 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1669;
              heapClock = ~ heapClock;
        end

       1669 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1002] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1670;
              heapClock = ~ heapClock;
        end

       1670 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[361] = localMem[1002];
              ip = 1671;
        end

       1671 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[5];
              heapArray  = localMem[361];
              heapIndex  = localMem[359];
              ip = 1672;
              heapClock = ~ heapClock;
        end

       1672 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1673;
              heapClock = ~ heapClock;
        end

       1673 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1003] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1674;
              heapClock = ~ heapClock;
        end

       1674 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1004] = localMem[1003] + 1;
              ip = 1675;
        end

       1675 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[355];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1004];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1676;
              heapClock = ~ heapClock;
        end

       1676 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 1690;
        end

       1677 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1678;
        end

       1678 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1679;
              heapClock = ~ heapClock;
        end

       1679 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1005] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1680;
              heapClock = ~ heapClock;
        end

       1680 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[362] = localMem[1005];
              ip = 1681;
        end

       1681 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[3];
              heapArray  = localMem[362];
              heapIndex  = localMem[357];
              ip = 1682;
              heapClock = ~ heapClock;
        end

       1682 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1683;
              heapClock = ~ heapClock;
        end

       1683 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1006] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1684;
              heapClock = ~ heapClock;
        end

       1684 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[363] = localMem[1006];
              ip = 1685;
        end

       1685 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[5];
              heapArray  = localMem[363];
              heapIndex  = localMem[357];
              ip = 1686;
              heapClock = ~ heapClock;
        end

       1686 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1687;
              heapClock = ~ heapClock;
        end

       1687 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1007] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1688;
              heapClock = ~ heapClock;
        end

       1688 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1008] = localMem[1007] + 1;
              ip = 1689;
        end

       1689 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[355];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1008];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1690;
              heapClock = ~ heapClock;
        end

       1690 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1691;
        end

       1691 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1692;
              heapClock = ~ heapClock;
        end

       1692 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1009] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1693;
              heapClock = ~ heapClock;
        end

       1693 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1010] = localMem[1009] + 1;
              ip = 1694;
        end

       1694 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[0];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1010];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1695;
              heapClock = ~ heapClock;
        end

       1695 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1696;
        end

       1696 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1697;
              heapClock = ~ heapClock;
        end

       1697 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1011] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1698;
              heapClock = ~ heapClock;
        end

       1698 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[365] = localMem[1011];
              ip = 1699;
        end

       1699 :
        begin                                                                   // jLt
          //$display("AAAA %4d %4d jLt", steps, ip);
              ip = localMem[365] <  3 ? 2159 : 1700;
        end

       1700 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1701;
              heapClock = ~ heapClock;
        end

       1701 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1012] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1702;
              heapClock = ~ heapClock;
        end

       1702 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[366] = localMem[1012];
              ip = 1703;
        end

       1703 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1704;
              heapClock = ~ heapClock;
        end

       1704 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1013] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1705;
              heapClock = ~ heapClock;
        end

       1705 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[367] = localMem[1013];
              ip = 1706;
        end

       1706 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[367] == 0 ? 1910 : 1707;
        end

       1707 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1708;
              heapClock = ~ heapClock;
        end

       1708 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[368] = heapOut;
              ip = 1709;
        end

       1709 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1014] = 1;
              ip = 1710;
        end

       1710 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1014];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1711;
              heapClock = ~ heapClock;
        end

       1711 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1015] = 0;
              ip = 1712;
        end

       1712 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1015];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1713;
              heapClock = ~ heapClock;
        end

       1713 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1714;
              heapClock = ~ heapClock;
        end

       1714 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[369] = heapOut;
              ip = 1715;
        end

       1715 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1016] = localMem[369];
              ip = 1716;
        end

       1716 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 4;                                                // Index of element to write to
              heapIn      = localMem[1016];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1717;
              heapClock = ~ heapClock;
        end

       1717 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 1718;
              heapClock = ~ heapClock;
        end

       1718 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[370] = heapOut;
              ip = 1719;
        end

       1719 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1017] = localMem[370];
              ip = 1720;
        end

       1720 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 5;                                                // Index of element to write to
              heapIn      = localMem[1017];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1721;
              heapClock = ~ heapClock;
        end

       1721 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1018] = 0;
              ip = 1722;
        end

       1722 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 6;                                                // Index of element to write to
              heapIn      = localMem[1018];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1723;
              heapClock = ~ heapClock;
        end

       1723 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1019] = localMem[366];
              ip = 1724;
        end

       1724 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 3;                                                // Index of element to write to
              heapIn      = localMem[1019];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1725;
              heapClock = ~ heapClock;
        end

       1725 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[366];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1726;
              heapClock = ~ heapClock;
        end

       1726 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1020] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1727;
              heapClock = ~ heapClock;
        end

       1727 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1021] = localMem[1020] + 1;
              ip = 1728;
        end

       1728 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[366];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1021];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1729;
              heapClock = ~ heapClock;
        end

       1729 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[366];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1730;
              heapClock = ~ heapClock;
        end

       1730 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1022] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1731;
              heapClock = ~ heapClock;
        end

       1731 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1023] = localMem[1022];
              ip = 1732;
        end

       1732 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1023];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1733;
              heapClock = ~ heapClock;
        end

       1733 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1734;
              heapClock = ~ heapClock;
        end

       1734 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1024] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1735;
              heapClock = ~ heapClock;
        end

       1735 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[371] = !localMem[1024];
              ip = 1736;
        end

       1736 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[371] != 0 ? 1791 : 1737;
        end

       1737 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1737");
        end

       1738 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1738");
        end

       1739 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1739");
        end

       1740 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1740");
        end

       1741 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1741");
        end

       1742 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1742");
        end

       1743 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1743");
        end

       1744 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1744");
        end

       1745 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1745");
        end

       1746 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1746");
        end

       1747 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1747");
        end

       1748 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1748");
        end

       1749 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1749");
        end

       1750 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1750");
        end

       1751 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1751");
        end

       1752 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1752");
        end

       1753 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1753");
        end

       1754 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1754");
        end

       1755 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1755");
        end

       1756 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1756");
        end

       1757 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1757");
        end

       1758 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1758");
        end

       1759 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1759");
        end

       1760 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1760");
        end

       1761 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1761");
        end

       1762 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1762");
        end

       1763 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1763");
        end

       1764 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1764");
        end

       1765 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1765");
        end

       1766 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1766");
        end

       1767 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1767");
        end

       1768 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1768");
        end

       1769 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1769");
        end

       1770 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1770");
        end

       1771 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1771");
        end

       1772 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1772");
        end

       1773 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1773");
        end

       1774 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1774");
        end

       1775 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1775");
        end

       1776 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  1776");
        end

       1777 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1777");
        end

       1778 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1778");
        end

       1779 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1779");
        end

       1780 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1780");
        end

       1781 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1781");
        end

       1782 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1782");
        end

       1783 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1783");
        end

       1784 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1784");
        end

       1785 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1785");
        end

       1786 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1786");
        end

       1787 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1787");
        end

       1788 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1788");
        end

       1789 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  1789");
        end

       1790 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1790");
        end

       1791 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1792;
        end

       1792 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1793;
              heapClock = ~ heapClock;
        end

       1793 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1037] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1794;
              heapClock = ~ heapClock;
        end

       1794 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[386] = localMem[1037];
              ip = 1795;
        end

       1795 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[368];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1796;
              heapClock = ~ heapClock;
        end

       1796 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1038] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1797;
              heapClock = ~ heapClock;
        end

       1797 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[387] = localMem[1038];
              ip = 1798;
        end

       1798 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[386];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1799;
              heapClock = ~ heapClock;
        end

       1799 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[387];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1800;
              heapClock = ~ heapClock;
        end

       1800 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1801;
              heapClock = ~ heapClock;
        end

       1801 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1039] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1802;
              heapClock = ~ heapClock;
        end

       1802 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[388] = localMem[1039];
              ip = 1803;
        end

       1803 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[368];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1804;
              heapClock = ~ heapClock;
        end

       1804 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1040] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1805;
              heapClock = ~ heapClock;
        end

       1805 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[389] = localMem[1040];
              ip = 1806;
        end

       1806 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[388];                                                 // Array to write to
              heapIndex  = 2;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 1807;
              heapClock = ~ heapClock;
        end

       1807 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[389];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 1;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 1808;
              heapClock = ~ heapClock;
        end

       1808 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1809;
        end

       1809 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1041] = 1;
              ip = 1810;
        end

       1810 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[355];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1041];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1811;
              heapClock = ~ heapClock;
        end

       1811 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1042] = localMem[367];
              ip = 1812;
        end

       1812 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[368];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1042];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1813;
              heapClock = ~ heapClock;
        end

       1813 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1814;
              heapClock = ~ heapClock;
        end

       1814 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1043] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1815;
              heapClock = ~ heapClock;
        end

       1815 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[390] = localMem[1043];
              ip = 1816;
        end

       1816 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1817;
              heapClock = ~ heapClock;
        end

       1817 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1044] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1818;
              heapClock = ~ heapClock;
        end

       1818 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[391] = localMem[1044];
              ip = 1819;
        end

       1819 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[391];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[390];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1820;
              heapClock = ~ heapClock;
        end

       1820 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1045] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1821;
              heapClock = ~ heapClock;
        end

       1821 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[392] = localMem[1045];
              ip = 1822;
        end

       1822 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[392] != localMem[355] ? 1863 : 1823;
        end

       1823 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1824;
              heapClock = ~ heapClock;
        end

       1824 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1046] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1825;
              heapClock = ~ heapClock;
        end

       1825 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[393] = localMem[1046];
              ip = 1826;
        end

       1826 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[393];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1827;
              heapClock = ~ heapClock;
        end

       1827 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1047] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1828;
              heapClock = ~ heapClock;
        end

       1828 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[394] = localMem[1047];
              ip = 1829;
        end

       1829 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1830;
              heapClock = ~ heapClock;
        end

       1830 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1048] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1831;
              heapClock = ~ heapClock;
        end

       1831 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[395] = localMem[1048];
              ip = 1832;
        end

       1832 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1049] = localMem[394];
              ip = 1833;
        end

       1833 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[395];                                                // Array to write to
              heapIndex   = localMem[390];                                                // Index of element to write to
              heapIn      = localMem[1049];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1834;
              heapClock = ~ heapClock;
        end

       1834 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1835;
              heapClock = ~ heapClock;
        end

       1835 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1050] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1836;
              heapClock = ~ heapClock;
        end

       1836 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[396] = localMem[1050];
              ip = 1837;
        end

       1837 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[396];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1838;
              heapClock = ~ heapClock;
        end

       1838 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1051] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1839;
              heapClock = ~ heapClock;
        end

       1839 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[397] = localMem[1051];
              ip = 1840;
        end

       1840 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1841;
              heapClock = ~ heapClock;
        end

       1841 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1052] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1842;
              heapClock = ~ heapClock;
        end

       1842 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[398] = localMem[1052];
              ip = 1843;
        end

       1843 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1053] = localMem[397];
              ip = 1844;
        end

       1844 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[398];                                                // Array to write to
              heapIndex   = localMem[390];                                                // Index of element to write to
              heapIn      = localMem[1053];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1845;
              heapClock = ~ heapClock;
        end

       1845 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1846;
              heapClock = ~ heapClock;
        end

       1846 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1054] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1847;
              heapClock = ~ heapClock;
        end

       1847 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[399] = localMem[1054];
              ip = 1848;
        end

       1848 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[399];
              ip = 1849;
              heapClock = ~ heapClock;
        end

       1849 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1850;
              heapClock = ~ heapClock;
        end

       1850 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1055] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1851;
              heapClock = ~ heapClock;
        end

       1851 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[400] = localMem[1055];
              ip = 1852;
        end

       1852 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[400];
              ip = 1853;
              heapClock = ~ heapClock;
        end

       1853 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[401] = localMem[390] + 1;
              ip = 1854;
        end

       1854 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1056] = localMem[401];
              ip = 1855;
        end

       1855 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[367];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1056];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1856;
              heapClock = ~ heapClock;
        end

       1856 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1857;
              heapClock = ~ heapClock;
        end

       1857 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1057] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1858;
              heapClock = ~ heapClock;
        end

       1858 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[402] = localMem[1057];
              ip = 1859;
        end

       1859 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1058] = localMem[368];
              ip = 1860;
        end

       1860 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[402];                                                // Array to write to
              heapIndex   = localMem[401];                                                // Index of element to write to
              heapIn      = localMem[1058];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1861;
              heapClock = ~ heapClock;
        end

       1861 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2156;
        end

       1862 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  1862");
        end

       1863 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 1864;
        end

       1864 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
            ip = 1865;
        end

       1865 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1866;
              heapClock = ~ heapClock;
        end

       1866 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1059] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1867;
              heapClock = ~ heapClock;
        end

       1867 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[403] = localMem[1059];
              ip = 1868;
        end

       1868 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[355];
              heapAction = `Index;
              heapArray  = localMem[403];
              ip = 1869;
              heapClock = ~ heapClock;
        end

       1869 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[404] = heapOut;
              ip = 1870;
        end

       1870 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[404] = localMem[404] - 1;
              ip = 1871;
        end

       1871 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1872;
              heapClock = ~ heapClock;
        end

       1872 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1060] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1873;
              heapClock = ~ heapClock;
        end

       1873 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[405] = localMem[1060];
              ip = 1874;
        end

       1874 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[405];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1875;
              heapClock = ~ heapClock;
        end

       1875 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1061] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1876;
              heapClock = ~ heapClock;
        end

       1876 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[406] = localMem[1061];
              ip = 1877;
        end

       1877 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1878;
              heapClock = ~ heapClock;
        end

       1878 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1062] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1879;
              heapClock = ~ heapClock;
        end

       1879 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[407] = localMem[1062];
              ip = 1880;
        end

       1880 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[407];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1881;
              heapClock = ~ heapClock;
        end

       1881 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1063] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1882;
              heapClock = ~ heapClock;
        end

       1882 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[408] = localMem[1063];
              ip = 1883;
        end

       1883 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1884;
              heapClock = ~ heapClock;
        end

       1884 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1064] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1885;
              heapClock = ~ heapClock;
        end

       1885 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[409] = localMem[1064];
              ip = 1886;
        end

       1886 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[409];
              ip = 1887;
              heapClock = ~ heapClock;
        end

       1887 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[355];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1888;
              heapClock = ~ heapClock;
        end

       1888 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1065] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1889;
              heapClock = ~ heapClock;
        end

       1889 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[410] = localMem[1065];
              ip = 1890;
        end

       1890 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
              heapAction = `Resize;
              heapIn     = 1;
              heapArray  = localMem[410];
              ip = 1891;
              heapClock = ~ heapClock;
        end

       1891 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1892;
              heapClock = ~ heapClock;
        end

       1892 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1066] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1893;
              heapClock = ~ heapClock;
        end

       1893 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[411] = localMem[1066];
              ip = 1894;
        end

       1894 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[406];
              heapArray  = localMem[411];
              heapIndex  = localMem[404];
              ip = 1895;
              heapClock = ~ heapClock;
        end

       1895 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1896;
              heapClock = ~ heapClock;
        end

       1896 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1067] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1897;
              heapClock = ~ heapClock;
        end

       1897 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[412] = localMem[1067];
              ip = 1898;
        end

       1898 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[408];
              heapArray  = localMem[412];
              heapIndex  = localMem[404];
              ip = 1899;
              heapClock = ~ heapClock;
        end

       1899 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1900;
              heapClock = ~ heapClock;
        end

       1900 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1068] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1901;
              heapClock = ~ heapClock;
        end

       1901 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[413] = localMem[1068];
              ip = 1902;
        end

       1902 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[414] = localMem[404] + 1;
              ip = 1903;
        end

       1903 :
        begin                                                                   // shiftUp
          //$display("AAAA %4d %4d shiftUp", steps, ip);
              heapAction = `Up;
              heapIn     = localMem[368];
              heapArray  = localMem[413];
              heapIndex  = localMem[414];
              ip = 1904;
              heapClock = ~ heapClock;
        end

       1904 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[367];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 1905;
              heapClock = ~ heapClock;
        end

       1905 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1069] = heapOut;                                                     // Data retrieved from heap memory
              ip = 1906;
              heapClock = ~ heapClock;
        end

       1906 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[1070] = localMem[1069] + 1;
              ip = 1907;
        end

       1907 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[367];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1070];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 1908;
              heapClock = ~ heapClock;
        end

       1908 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2156;
        end

       1909 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1909");
        end

       1910 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  1910");
        end

       1911 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1911");
        end

       1912 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1912");
        end

       1913 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1913");
        end

       1914 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1914");
        end

       1915 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1915");
        end

       1916 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1916");
        end

       1917 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1917");
        end

       1918 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1918");
        end

       1919 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1919");
        end

       1920 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1920");
        end

       1921 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1921");
        end

       1922 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1922");
        end

       1923 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1923");
        end

       1924 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1924");
        end

       1925 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1925");
        end

       1926 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1926");
        end

       1927 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1927");
        end

       1928 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1928");
        end

       1929 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1929");
        end

       1930 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1930");
        end

       1931 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1931");
        end

       1932 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1932");
        end

       1933 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1933");
        end

       1934 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1934");
        end

       1935 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1935");
        end

       1936 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1936");
        end

       1937 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1937");
        end

       1938 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1938");
        end

       1939 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1939");
        end

       1940 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1940");
        end

       1941 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1941");
        end

       1942 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1942");
        end

       1943 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1943");
        end

       1944 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1944");
        end

       1945 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1945");
        end

       1946 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1946");
        end

       1947 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1947");
        end

       1948 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1948");
        end

       1949 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1949");
        end

       1950 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1950");
        end

       1951 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1951");
        end

       1952 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1952");
        end

       1953 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1953");
        end

       1954 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1954");
        end

       1955 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1955");
        end

       1956 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1956");
        end

       1957 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1957");
        end

       1958 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1958");
        end

       1959 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1959");
        end

       1960 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1960");
        end

       1961 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1961");
        end

       1962 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1962");
        end

       1963 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1963");
        end

       1964 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1964");
        end

       1965 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
          // $display("Should not be executed  1965");
        end

       1966 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
          // $display("Should not be executed  1966");
        end

       1967 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1967");
        end

       1968 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1968");
        end

       1969 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1969");
        end

       1970 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1970");
        end

       1971 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  1971");
        end

       1972 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  1972");
        end

       1973 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1973");
        end

       1974 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  1974");
        end

       1975 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1975");
        end

       1976 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1976");
        end

       1977 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1977");
        end

       1978 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1978");
        end

       1979 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1979");
        end

       1980 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1980");
        end

       1981 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1981");
        end

       1982 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1982");
        end

       1983 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1983");
        end

       1984 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1984");
        end

       1985 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1985");
        end

       1986 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1986");
        end

       1987 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1987");
        end

       1988 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1988");
        end

       1989 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1989");
        end

       1990 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1990");
        end

       1991 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1991");
        end

       1992 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1992");
        end

       1993 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1993");
        end

       1994 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  1994");
        end

       1995 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  1995");
        end

       1996 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  1996");
        end

       1997 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  1997");
        end

       1998 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  1998");
        end

       1999 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  1999");
        end

       2000 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2000");
        end

       2001 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2001");
        end

       2002 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2002");
        end

       2003 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2003");
        end

       2004 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2004");
        end

       2005 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2005");
        end

       2006 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2006");
        end

       2007 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2007");
        end

       2008 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2008");
        end

       2009 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2009");
        end

       2010 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2010");
        end

       2011 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2011");
        end

       2012 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2012");
        end

       2013 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2013");
        end

       2014 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2014");
        end

       2015 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2015");
        end

       2016 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2016");
        end

       2017 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2017");
        end

       2018 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2018");
        end

       2019 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2019");
        end

       2020 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2020");
        end

       2021 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2021");
        end

       2022 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2022");
        end

       2023 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2023");
        end

       2024 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2024");
        end

       2025 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2025");
        end

       2026 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2026");
        end

       2027 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2027");
        end

       2028 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2028");
        end

       2029 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2029");
        end

       2030 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2030");
        end

       2031 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2031");
        end

       2032 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2032");
        end

       2033 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2033");
        end

       2034 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2034");
        end

       2035 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2035");
        end

       2036 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2036");
        end

       2037 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2037");
        end

       2038 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2038");
        end

       2039 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2039");
        end

       2040 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2040");
        end

       2041 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2041");
        end

       2042 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2042");
        end

       2043 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2043");
        end

       2044 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2044");
        end

       2045 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2045");
        end

       2046 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2046");
        end

       2047 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2047");
        end

       2048 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2048");
        end

       2049 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2049");
        end

       2050 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2050");
        end

       2051 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2051");
        end

       2052 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2052");
        end

       2053 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2053");
        end

       2054 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2054");
        end

       2055 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
          // $display("Should not be executed  2055");
        end

       2056 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2056");
        end

       2057 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2057");
        end

       2058 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2058");
        end

       2059 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2059");
        end

       2060 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2060");
        end

       2061 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2061");
        end

       2062 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
          // $display("Should not be executed  2062");
        end

       2063 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2063");
        end

       2064 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2064");
        end

       2065 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2065");
        end

       2066 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2066");
        end

       2067 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
          // $display("Should not be executed  2067");
        end

       2068 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
          // $display("Should not be executed  2068");
        end

       2069 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2069");
        end

       2070 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2070");
        end

       2071 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2071");
        end

       2072 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2072");
        end

       2073 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2073");
        end

       2074 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2074");
        end

       2075 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2075");
        end

       2076 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2076");
        end

       2077 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2077");
        end

       2078 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2078");
        end

       2079 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2079");
        end

       2080 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2080");
        end

       2081 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2081");
        end

       2082 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2082");
        end

       2083 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2083");
        end

       2084 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2084");
        end

       2085 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2085");
        end

       2086 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2086");
        end

       2087 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2087");
        end

       2088 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2088");
        end

       2089 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2089");
        end

       2090 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2090");
        end

       2091 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2091");
        end

       2092 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2092");
        end

       2093 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2093");
        end

       2094 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2094");
        end

       2095 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2095");
        end

       2096 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2096");
        end

       2097 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2097");
        end

       2098 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2098");
        end

       2099 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2099");
        end

       2100 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2100");
        end

       2101 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
          // $display("Should not be executed  2101");
        end

       2102 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
          // $display("Should not be executed  2102");
        end

       2103 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2103");
        end

       2104 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2104");
        end

       2105 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2105");
        end

       2106 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2106");
        end

       2107 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2107");
        end

       2108 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2108");
        end

       2109 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2109");
        end

       2110 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2110");
        end

       2111 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2111");
        end

       2112 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2112");
        end

       2113 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2113");
        end

       2114 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2114");
        end

       2115 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2115");
        end

       2116 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2116");
        end

       2117 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2117");
        end

       2118 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2118");
        end

       2119 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2119");
        end

       2120 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2120");
        end

       2121 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2121");
        end

       2122 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2122");
        end

       2123 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2123");
        end

       2124 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2124");
        end

       2125 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2125");
        end

       2126 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2126");
        end

       2127 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2127");
        end

       2128 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2128");
        end

       2129 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2129");
        end

       2130 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2130");
        end

       2131 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2131");
        end

       2132 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2132");
        end

       2133 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2133");
        end

       2134 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2134");
        end

       2135 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2135");
        end

       2136 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2136");
        end

       2137 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2137");
        end

       2138 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2138");
        end

       2139 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2139");
        end

       2140 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2140");
        end

       2141 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2141");
        end

       2142 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2142");
        end

       2143 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2143");
        end

       2144 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2144");
        end

       2145 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2145");
        end

       2146 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2146");
        end

       2147 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2147");
        end

       2148 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2148");
        end

       2149 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2149");
        end

       2150 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
          // $display("Should not be executed  2150");
        end

       2151 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
          // $display("Should not be executed  2151");
        end

       2152 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2152");
        end

       2153 :
        begin                                                                   // resize
          //$display("AAAA %4d %4d resize", steps, ip);
          // $display("Should not be executed  2153");
        end

       2154 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2154");
        end

       2155 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2155");
        end

       2156 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2157;
        end

       2157 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[364] = 1;
              ip = 2158;
        end

       2158 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2161;
        end

       2159 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2160;
        end

       2160 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[364] = 0;
              ip = 2161;
        end

       2161 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2162;
        end

       2162 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2163;
        end

       2163 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2164;
        end

       2164 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2165;
        end

       2165 :
        begin                                                                   // tally
          //$display("AAAA %4d %4d tally", steps, ip);
            ip = 2166;
        end

       2166 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2167;
        end

       2167 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 14;
        end

       2168 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2169;
        end

       2169 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[468] = 1;
              ip = 2170;
        end

       2170 :
        begin                                                                   // shiftLeft
          //$display("AAAA %4d %4d shiftLeft", steps, ip);
              localMem[468] = localMem[468] << 31;
              ip = 2171;
        end

       2171 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2172;
              heapClock = ~ heapClock;
        end

       2172 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1141] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2173;
              heapClock = ~ heapClock;
        end

       2173 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[469] = localMem[1141];
              ip = 2174;
        end

       2174 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2175;
              heapClock = ~ heapClock;
        end

       2175 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[470] = heapOut;
              ip = 2176;
        end

       2176 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2177;
              heapClock = ~ heapClock;
        end

       2177 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[471] = heapOut;
              ip = 2178;
        end

       2178 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[469] != 0 ? 2186 : 2179;
        end

       2179 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2179");
        end

       2180 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2180");
        end

       2181 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2181");
        end

       2182 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2182");
        end

       2183 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2183");
        end

       2184 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2184");
        end

       2185 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2185");
        end

       2186 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2187;
        end

       2187 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2188;
        end

       2188 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[472] = 0;
              ip = 2189;
        end

       2189 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2190;
        end

       2190 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[472] >= 99 ? 2205 : 2191;
        end

       2191 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[469];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2192;
              heapClock = ~ heapClock;
        end

       2192 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1145] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2193;
              heapClock = ~ heapClock;
        end

       2193 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[473] = !localMem[1145];
              ip = 2194;
        end

       2194 :
        begin                                                                   // jTrue
          //$display("AAAA %4d %4d jTrue", steps, ip);
              ip = localMem[473] != 0 ? 2205 : 2195;
        end

       2195 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[469];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2196;
              heapClock = ~ heapClock;
        end

       2196 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1146] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2197;
              heapClock = ~ heapClock;
        end

       2197 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[474] = localMem[1146];
              ip = 2198;
        end

       2198 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[474];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2199;
              heapClock = ~ heapClock;
        end

       2199 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1147] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2200;
              heapClock = ~ heapClock;
        end

       2200 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[475] = localMem[1147];
              ip = 2201;
        end

       2201 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[469] = localMem[475];
              ip = 2202;
        end

       2202 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2203;
        end

       2203 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[472] = localMem[472] + 1;
              ip = 2204;
        end

       2204 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2189;
        end

       2205 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2206;
        end

       2206 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1148] = localMem[469];
              ip = 2207;
        end

       2207 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1148];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2208;
              heapClock = ~ heapClock;
        end

       2208 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1149] = 1;
              ip = 2209;
        end

       2209 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1149];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2210;
              heapClock = ~ heapClock;
        end

       2210 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1150] = 0;
              ip = 2211;
        end

       2211 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1150];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2212;
              heapClock = ~ heapClock;
        end

       2212 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2213;
        end

       2213 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2214;
        end

       2214 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[470];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2215;
              heapClock = ~ heapClock;
        end

       2215 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1151] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2216;
              heapClock = ~ heapClock;
        end

       2216 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[476] = localMem[1151];
              ip = 2217;
        end

       2217 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[476] == 3 ? 2457 : 2218;
        end

       2218 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[470];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 2219;
              heapClock = ~ heapClock;
        end

       2219 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[471];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 3;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 2220;
              heapClock = ~ heapClock;
        end

       2220 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[471];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2221;
              heapClock = ~ heapClock;
        end

       2221 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1152] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2222;
              heapClock = ~ heapClock;
        end

       2222 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[477] = localMem[1152];
              ip = 2223;
        end

       2223 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[471];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2224;
              heapClock = ~ heapClock;
        end

       2224 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1153] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2225;
              heapClock = ~ heapClock;
        end

       2225 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[478] = localMem[1153];
              ip = 2226;
        end

       2226 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[477];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2227;
              heapClock = ~ heapClock;
        end

       2227 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1154] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2228;
              heapClock = ~ heapClock;
        end

       2228 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[479] = localMem[1154];
              ip = 2229;
        end

       2229 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[479];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[478];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2230;
              heapClock = ~ heapClock;
        end

       2230 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1155] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2231;
              heapClock = ~ heapClock;
        end

       2231 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[480] = localMem[1155];
              ip = 2232;
        end

       2232 :
        begin                                                                   // out
          //$display("AAAA %4d %4d out", steps, ip);
              outMem[outMemPos] = localMem[480];
              outMemPos = outMemPos + 1;
              ip = 2233;
        end

       2233 :
        begin                                                                   // tally
          //$display("AAAA %4d %4d tally", steps, ip);
            ip = 2234;
        end

       2234 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2235;
        end

       2235 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2236;
              heapClock = ~ heapClock;
        end

       2236 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1156] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2237;
              heapClock = ~ heapClock;
        end

       2237 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = localMem[1156];
              ip = 2238;
        end

       2238 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[481] != 0 ? 2246 : 2239;
        end

       2239 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2239");
        end

       2240 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2240");
        end

       2241 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2241");
        end

       2242 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2242");
        end

       2243 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2243");
        end

       2244 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2244");
        end

       2245 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2245");
        end

       2246 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2247;
        end

       2247 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2248;
        end

       2248 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[482] = 0;
              ip = 2249;
        end

       2249 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2250;
        end

       2250 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[482] >= 99 ? 2317 : 2251;
        end

       2251 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2252;
              heapClock = ~ heapClock;
        end

       2252 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1160] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2253;
              heapClock = ~ heapClock;
        end

       2253 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[483] = localMem[1160] - 1;
              ip = 2254;
        end

       2254 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 4;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2255;
              heapClock = ~ heapClock;
        end

       2255 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1161] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2256;
              heapClock = ~ heapClock;
        end

       2256 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[484] = localMem[1161];
              ip = 2257;
        end

       2257 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[484];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[483];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2258;
              heapClock = ~ heapClock;
        end

       2258 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1162] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2259;
              heapClock = ~ heapClock;
        end

       2259 :
        begin                                                                   // jLe
          //$display("AAAA %4d %4d jLe", steps, ip);
              ip = localMem[480] <= localMem[1162] ? 2281 : 2260;
        end

       2260 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[485] = localMem[483] + 1;
              ip = 2261;
        end

       2261 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2262;
              heapClock = ~ heapClock;
        end

       2262 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1163] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2263;
              heapClock = ~ heapClock;
        end

       2263 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[486] = !localMem[1163];
              ip = 2264;
        end

       2264 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[486] == 0 ? 2272 : 2265;
        end

       2265 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2265");
        end

       2266 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2266");
        end

       2267 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2267");
        end

       2268 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2268");
        end

       2269 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2269");
        end

       2270 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2270");
        end

       2271 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2271");
        end

       2272 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2273;
        end

       2273 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2274;
              heapClock = ~ heapClock;
        end

       2274 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1167] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2275;
              heapClock = ~ heapClock;
        end

       2275 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[487] = localMem[1167];
              ip = 2276;
        end

       2276 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[487];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[485];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2277;
              heapClock = ~ heapClock;
        end

       2277 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1168] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2278;
              heapClock = ~ heapClock;
        end

       2278 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[488] = localMem[1168];
              ip = 2279;
        end

       2279 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = localMem[488];
              ip = 2280;
        end

       2280 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2314;
        end

       2281 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2282;
        end

       2282 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[480];
              heapAction = `Index;
              heapArray  = localMem[484];
              ip = 2283;
              heapClock = ~ heapClock;
        end

       2283 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[489] = heapOut;
              ip = 2284;
        end

       2284 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[489] == 0 ? 2292 : 2285;
        end

       2285 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1169] = localMem[481];
              ip = 2286;
        end

       2286 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1169];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2287;
              heapClock = ~ heapClock;
        end

       2287 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1170] = 1;
              ip = 2288;
        end

       2288 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1170];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2289;
              heapClock = ~ heapClock;
        end

       2289 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[1171] = localMem[489] - 1;
              ip = 2290;
        end

       2290 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[1];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1171];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2291;
              heapClock = ~ heapClock;
        end

       2291 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2321;
        end

       2292 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2293;
        end

       2293 :
        begin                                                                   // arrayCountLess
          //$display("AAAA %4d %4d arrayCountLess", steps, ip);
              heapIn     = localMem[480];
              heapAction = `Less;
              heapArray  = localMem[484];
              ip = 2294;
              heapClock = ~ heapClock;
        end

       2294 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[490] = heapOut;
              ip = 2295;
        end

       2295 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2296;
              heapClock = ~ heapClock;
        end

       2296 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1172] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2297;
              heapClock = ~ heapClock;
        end

       2297 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[491] = !localMem[1172];
              ip = 2298;
        end

       2298 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[491] == 0 ? 2306 : 2299;
        end

       2299 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2299");
        end

       2300 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2300");
        end

       2301 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2301");
        end

       2302 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2302");
        end

       2303 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2303");
        end

       2304 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2304");
        end

       2305 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2305");
        end

       2306 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2307;
        end

       2307 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[481];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2308;
              heapClock = ~ heapClock;
        end

       2308 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1176] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2309;
              heapClock = ~ heapClock;
        end

       2309 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[492] = localMem[1176];
              ip = 2310;
        end

       2310 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[492];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[490];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2311;
              heapClock = ~ heapClock;
        end

       2311 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1177] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2312;
              heapClock = ~ heapClock;
        end

       2312 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[493] = localMem[1177];
              ip = 2313;
        end

       2313 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[481] = localMem[493];
              ip = 2314;
        end

       2314 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2315;
        end

       2315 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[482] = localMem[482] + 1;
              ip = 2316;
        end

       2316 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2249;
        end

       2317 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2317");
        end

       2318 :
        begin                                                                   // assert
          //$display("AAAA %4d %4d assert", steps, ip);
          // $display("Should not be executed  2318");
        end

       2319 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2319");
        end

       2320 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2320");
        end

       2321 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2322;
        end

       2322 :
        begin                                                                   // tally
          //$display("AAAA %4d %4d tally", steps, ip);
            ip = 2323;
        end

       2323 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[1];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2324;
              heapClock = ~ heapClock;
        end

       2324 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1178] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2325;
              heapClock = ~ heapClock;
        end

       2325 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[494] = localMem[1178];
              ip = 2326;
        end

       2326 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[1];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2327;
              heapClock = ~ heapClock;
        end

       2327 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1179] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2328;
              heapClock = ~ heapClock;
        end

       2328 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[495] = localMem[1179];
              ip = 2329;
        end

       2329 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[494];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 5;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2330;
              heapClock = ~ heapClock;
        end

       2330 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1180] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2331;
              heapClock = ~ heapClock;
        end

       2331 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[496] = localMem[1180];
              ip = 2332;
        end

       2332 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[496];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[495];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2333;
              heapClock = ~ heapClock;
        end

       2333 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1181] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2334;
              heapClock = ~ heapClock;
        end

       2334 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[497] = localMem[1181];
              ip = 2335;
        end

       2335 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[498] = localMem[480] + localMem[480];
              ip = 2336;
        end

       2336 :
        begin                                                                   // assertEq
          //$display("AAAA %4d %4d assertEq", steps, ip);
            ip = 2337;
        end

       2337 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2338;
        end

       2338 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[470];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2339;
              heapClock = ~ heapClock;
        end

       2339 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1182] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2340;
              heapClock = ~ heapClock;
        end

       2340 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[499] = localMem[1182];
              ip = 2341;
        end

       2341 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2342;
              heapClock = ~ heapClock;
        end

       2342 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1183] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2343;
              heapClock = ~ heapClock;
        end

       2343 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[500] = !localMem[1183];
              ip = 2344;
        end

       2344 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[500] == 0 ? 2406 : 2345;
        end

       2345 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[470];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2346;
              heapClock = ~ heapClock;
        end

       2346 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1184] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2347;
              heapClock = ~ heapClock;
        end

       2347 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[501] = localMem[1184] + 1;
              ip = 2348;
        end

       2348 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2349;
              heapClock = ~ heapClock;
        end

       2349 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1185] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2350;
              heapClock = ~ heapClock;
        end

       2350 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[502] = localMem[1185];
              ip = 2351;
        end

       2351 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[501] >= localMem[502] ? 2359 : 2352;
        end

       2352 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1186] = localMem[499];
              ip = 2353;
        end

       2353 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1186];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2354;
              heapClock = ~ heapClock;
        end

       2354 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1187] = 1;
              ip = 2355;
        end

       2355 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1187];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2356;
              heapClock = ~ heapClock;
        end

       2356 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1188] = localMem[501];
              ip = 2357;
        end

       2357 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1188];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2358;
              heapClock = ~ heapClock;
        end

       2358 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2453;
        end

       2359 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2360;
        end

       2360 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2361;
              heapClock = ~ heapClock;
        end

       2361 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1189] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2362;
              heapClock = ~ heapClock;
        end

       2362 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[503] = localMem[1189];
              ip = 2363;
        end

       2363 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[503] == 0 ? 2398 : 2364;
        end

       2364 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2365;
        end

       2365 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[504] = 0;
              ip = 2366;
        end

       2366 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2367;
        end

       2367 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[504] >= 99 ? 2397 : 2368;
        end

       2368 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[503];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2369;
              heapClock = ~ heapClock;
        end

       2369 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1190] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2370;
              heapClock = ~ heapClock;
        end

       2370 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[505] = localMem[1190];
              ip = 2371;
        end

       2371 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
            ip = 2372;
        end

       2372 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[503];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2373;
              heapClock = ~ heapClock;
        end

       2373 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1191] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2374;
              heapClock = ~ heapClock;
        end

       2374 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[506] = localMem[1191];
              ip = 2375;
        end

       2375 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[499];
              heapAction = `Index;
              heapArray  = localMem[506];
              ip = 2376;
              heapClock = ~ heapClock;
        end

       2376 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[507] = heapOut;
              ip = 2377;
        end

       2377 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[507] = localMem[507] - 1;
              ip = 2378;
        end

       2378 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[507] != localMem[505] ? 2385 : 2379;
        end

       2379 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[499] = localMem[503];
              ip = 2380;
        end

       2380 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2381;
              heapClock = ~ heapClock;
        end

       2381 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1192] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2382;
              heapClock = ~ heapClock;
        end

       2382 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[503] = localMem[1192];
              ip = 2383;
        end

       2383 :
        begin                                                                   // jFalse
          //$display("AAAA %4d %4d jFalse", steps, ip);
              ip = localMem[503] == 0 ? 2397 : 2384;
        end

       2384 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2393;
        end

       2385 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2386;
        end

       2386 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1193] = localMem[503];
              ip = 2387;
        end

       2387 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1193];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2388;
              heapClock = ~ heapClock;
        end

       2388 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1194] = 1;
              ip = 2389;
        end

       2389 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1194];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2390;
              heapClock = ~ heapClock;
        end

       2390 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1195] = localMem[507];
              ip = 2391;
        end

       2391 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1195];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2392;
              heapClock = ~ heapClock;
        end

       2392 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2453;
        end

       2393 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2394;
        end

       2394 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2395;
        end

       2395 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[504] = localMem[504] + 1;
              ip = 2396;
        end

       2396 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2366;
        end

       2397 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2398;
        end

       2398 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2399;
        end

       2399 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1196] = localMem[499];
              ip = 2400;
        end

       2400 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1196];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2401;
              heapClock = ~ heapClock;
        end

       2401 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1197] = 3;
              ip = 2402;
        end

       2402 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1197];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2403;
              heapClock = ~ heapClock;
        end

       2403 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1198] = 0;
              ip = 2404;
        end

       2404 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1198];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2405;
              heapClock = ~ heapClock;
        end

       2405 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2453;
        end

       2406 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2407;
        end

       2407 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[470];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2408;
              heapClock = ~ heapClock;
        end

       2408 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1199] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2409;
              heapClock = ~ heapClock;
        end

       2409 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[508] = localMem[1199] + 1;
              ip = 2410;
        end

       2410 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[499];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2411;
              heapClock = ~ heapClock;
        end

       2411 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1200] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2412;
              heapClock = ~ heapClock;
        end

       2412 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[509] = localMem[1200];
              ip = 2413;
        end

       2413 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[509];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[508];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2414;
              heapClock = ~ heapClock;
        end

       2414 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1201] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2415;
              heapClock = ~ heapClock;
        end

       2415 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[510] = localMem[1201];
              ip = 2416;
        end

       2416 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[510] != 0 ? 2424 : 2417;
        end

       2417 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2417");
        end

       2418 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2418");
        end

       2419 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2419");
        end

       2420 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2420");
        end

       2421 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2421");
        end

       2422 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2422");
        end

       2423 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2423");
        end

       2424 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2425;
        end

       2425 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2426;
        end

       2426 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[511] = 0;
              ip = 2427;
        end

       2427 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2428;
        end

       2428 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[511] >= 99 ? 2443 : 2429;
        end

       2429 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[510];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2430;
              heapClock = ~ heapClock;
        end

       2430 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1205] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2431;
              heapClock = ~ heapClock;
        end

       2431 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[512] = !localMem[1205];
              ip = 2432;
        end

       2432 :
        begin                                                                   // jTrue
          //$display("AAAA %4d %4d jTrue", steps, ip);
              ip = localMem[512] != 0 ? 2443 : 2433;
        end

       2433 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[510];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2434;
              heapClock = ~ heapClock;
        end

       2434 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1206] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2435;
              heapClock = ~ heapClock;
        end

       2435 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[513] = localMem[1206];
              ip = 2436;
        end

       2436 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[513];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2437;
              heapClock = ~ heapClock;
        end

       2437 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1207] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2438;
              heapClock = ~ heapClock;
        end

       2438 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[514] = localMem[1207];
              ip = 2439;
        end

       2439 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[510] = localMem[514];
              ip = 2440;
        end

       2440 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2441;
        end

       2441 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[511] = localMem[511] + 1;
              ip = 2442;
        end

       2442 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2427;
        end

       2443 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2444;
        end

       2444 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1208] = localMem[510];
              ip = 2445;
        end

       2445 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1208];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2446;
              heapClock = ~ heapClock;
        end

       2446 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1209] = 1;
              ip = 2447;
        end

       2447 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1209];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2448;
              heapClock = ~ heapClock;
        end

       2448 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1210] = 0;
              ip = 2449;
        end

       2449 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[470];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1210];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2450;
              heapClock = ~ heapClock;
        end

       2450 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2451;
        end

       2451 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2452;
        end

       2452 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2453;
        end

       2453 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2454;
        end

       2454 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2213;
        end

       2455 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2455");
        end

       2456 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2456");
        end

       2457 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2458;
        end

       2458 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[470];
              ip = 2459;
              heapClock = ~ heapClock;
        end

       2459 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[471];
              ip = 2460;
              heapClock = ~ heapClock;
        end

       2460 :
        begin                                                                   // tally
          //$display("AAAA %4d %4d tally", steps, ip);
            ip = 2461;
        end

       2461 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[515] = 1;
              ip = 2462;
        end

       2462 :
        begin                                                                   // shiftLeft
          //$display("AAAA %4d %4d shiftLeft", steps, ip);
              localMem[515] = localMem[515] << 31;
              ip = 2463;
        end

       2463 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[0];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 3;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2464;
              heapClock = ~ heapClock;
        end

       2464 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1211] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2465;
              heapClock = ~ heapClock;
        end

       2465 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[516] = localMem[1211];
              ip = 2466;
        end

       2466 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2467;
              heapClock = ~ heapClock;
        end

       2467 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[517] = heapOut;
              ip = 2468;
        end

       2468 :
        begin                                                                   // array
          //$display("AAAA %4d %4d array", steps, ip);
              heapAction = `Alloc;
              ip = 2469;
              heapClock = ~ heapClock;
        end

       2469 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[518] = heapOut;
              ip = 2470;
        end

       2470 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[516] != 0 ? 2478 : 2471;
        end

       2471 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2471");
        end

       2472 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2472");
        end

       2473 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2473");
        end

       2474 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2474");
        end

       2475 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2475");
        end

       2476 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2476");
        end

       2477 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2477");
        end

       2478 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2479;
        end

       2479 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2480;
        end

       2480 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[519] = 0;
              ip = 2481;
        end

       2481 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2482;
        end

       2482 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[519] >= 99 ? 2497 : 2483;
        end

       2483 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[516];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2484;
              heapClock = ~ heapClock;
        end

       2484 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1215] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2485;
              heapClock = ~ heapClock;
        end

       2485 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[520] = !localMem[1215];
              ip = 2486;
        end

       2486 :
        begin                                                                   // jTrue
          //$display("AAAA %4d %4d jTrue", steps, ip);
              ip = localMem[520] != 0 ? 2497 : 2487;
        end

       2487 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[516];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2488;
              heapClock = ~ heapClock;
        end

       2488 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1216] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2489;
              heapClock = ~ heapClock;
        end

       2489 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[521] = localMem[1216];
              ip = 2490;
        end

       2490 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[521];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2491;
              heapClock = ~ heapClock;
        end

       2491 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1217] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2492;
              heapClock = ~ heapClock;
        end

       2492 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[522] = localMem[1217];
              ip = 2493;
        end

       2493 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[516] = localMem[522];
              ip = 2494;
        end

       2494 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2495;
        end

       2495 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[519] = localMem[519] + 1;
              ip = 2496;
        end

       2496 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2481;
        end

       2497 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2498;
        end

       2498 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1218] = localMem[516];
              ip = 2499;
        end

       2499 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1218];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2500;
              heapClock = ~ heapClock;
        end

       2500 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1219] = 1;
              ip = 2501;
        end

       2501 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1219];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2502;
              heapClock = ~ heapClock;
        end

       2502 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1220] = 0;
              ip = 2503;
        end

       2503 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1220];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2504;
              heapClock = ~ heapClock;
        end

       2504 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2505;
        end

       2505 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2506;
        end

       2506 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[517];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 1;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2507;
              heapClock = ~ heapClock;
        end

       2507 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1221] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2508;
              heapClock = ~ heapClock;
        end

       2508 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[523] = localMem[1221];
              ip = 2509;
        end

       2509 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[523] == 3 ? 2632 : 2510;
        end

       2510 :
        begin                                                                   // moveLong1
          //$display("AAAA %4d %4d moveLong1", steps, ip);
              heapArray  = localMem[517];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapAction = `Long1;                                          // Request a write
              ip = 2511;
              heapClock = ~ heapClock;
        end

       2511 :
        begin                                                                   // moveLong2
          //$display("AAAA %4d %4d moveLong2", steps, ip);
              heapArray  = localMem[518];                                                 // Array to write to
              heapIndex  = 0;                                                 // Index of element to write to
              heapIn     = 3;                                                  // Index of element to write to
              heapAction = `Long2;                                          // Request a write
              ip = 2512;
              heapClock = ~ heapClock;
        end

       2512 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2513;
        end

       2513 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[517];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2514;
              heapClock = ~ heapClock;
        end

       2514 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1222] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2515;
              heapClock = ~ heapClock;
        end

       2515 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[524] = localMem[1222];
              ip = 2516;
        end

       2516 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[524];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2517;
              heapClock = ~ heapClock;
        end

       2517 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1223] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2518;
              heapClock = ~ heapClock;
        end

       2518 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[525] = !localMem[1223];
              ip = 2519;
        end

       2519 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[525] == 0 ? 2581 : 2520;
        end

       2520 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[517];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2521;
              heapClock = ~ heapClock;
        end

       2521 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1224] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2522;
              heapClock = ~ heapClock;
        end

       2522 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[526] = localMem[1224] + 1;
              ip = 2523;
        end

       2523 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[524];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2524;
              heapClock = ~ heapClock;
        end

       2524 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1225] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2525;
              heapClock = ~ heapClock;
        end

       2525 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[527] = localMem[1225];
              ip = 2526;
        end

       2526 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[526] >= localMem[527] ? 2534 : 2527;
        end

       2527 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1226] = localMem[524];
              ip = 2528;
        end

       2528 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1226];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2529;
              heapClock = ~ heapClock;
        end

       2529 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1227] = 1;
              ip = 2530;
        end

       2530 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1227];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2531;
              heapClock = ~ heapClock;
        end

       2531 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1228] = localMem[526];
              ip = 2532;
        end

       2532 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1228];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2533;
              heapClock = ~ heapClock;
        end

       2533 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2628;
        end

       2534 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2535;
        end

       2535 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[524];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2536;
              heapClock = ~ heapClock;
        end

       2536 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1229] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2537;
              heapClock = ~ heapClock;
        end

       2537 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[528] = localMem[1229];
              ip = 2538;
        end

       2538 :
        begin                                                                   // jEq
          //$display("AAAA %4d %4d jEq", steps, ip);
              ip = localMem[528] == 0 ? 2573 : 2539;
        end

       2539 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2540;
        end

       2540 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[529] = 0;
              ip = 2541;
        end

       2541 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2542;
        end

       2542 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[529] >= 99 ? 2572 : 2543;
        end

       2543 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[528];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2544;
              heapClock = ~ heapClock;
        end

       2544 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1230] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2545;
              heapClock = ~ heapClock;
        end

       2545 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[530] = localMem[1230];
              ip = 2546;
        end

       2546 :
        begin                                                                   // assertNe
          //$display("AAAA %4d %4d assertNe", steps, ip);
            ip = 2547;
        end

       2547 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[528];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2548;
              heapClock = ~ heapClock;
        end

       2548 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1231] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2549;
              heapClock = ~ heapClock;
        end

       2549 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[531] = localMem[1231];
              ip = 2550;
        end

       2550 :
        begin                                                                   // arrayIndex
          //$display("AAAA %4d %4d arrayIndex", steps, ip);
              heapIn     = localMem[524];
              heapAction = `Index;
              heapArray  = localMem[531];
              ip = 2551;
              heapClock = ~ heapClock;
        end

       2551 :
        begin                                                                   // movHeapOut
          //$display("AAAA %4d %4d movHeapOut", steps, ip);
              localMem[532] = heapOut;
              ip = 2552;
        end

       2552 :
        begin                                                                   // subtract
          //$display("AAAA %4d %4d subtract", steps, ip);
              localMem[532] = localMem[532] - 1;
              ip = 2553;
        end

       2553 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[532] != localMem[530] ? 2560 : 2554;
        end

       2554 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[524] = localMem[528];
              ip = 2555;
        end

       2555 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[524];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2556;
              heapClock = ~ heapClock;
        end

       2556 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1232] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2557;
              heapClock = ~ heapClock;
        end

       2557 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[528] = localMem[1232];
              ip = 2558;
        end

       2558 :
        begin                                                                   // jFalse
          //$display("AAAA %4d %4d jFalse", steps, ip);
              ip = localMem[528] == 0 ? 2572 : 2559;
        end

       2559 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2568;
        end

       2560 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2561;
        end

       2561 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1233] = localMem[528];
              ip = 2562;
        end

       2562 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1233];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2563;
              heapClock = ~ heapClock;
        end

       2563 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1234] = 1;
              ip = 2564;
        end

       2564 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1234];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2565;
              heapClock = ~ heapClock;
        end

       2565 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1235] = localMem[532];
              ip = 2566;
        end

       2566 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1235];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2567;
              heapClock = ~ heapClock;
        end

       2567 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2628;
        end

       2568 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2569;
        end

       2569 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2570;
        end

       2570 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[529] = localMem[529] + 1;
              ip = 2571;
        end

       2571 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2541;
        end

       2572 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2573;
        end

       2573 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2574;
        end

       2574 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1236] = localMem[524];
              ip = 2575;
        end

       2575 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1236];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2576;
              heapClock = ~ heapClock;
        end

       2576 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1237] = 3;
              ip = 2577;
        end

       2577 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1237];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2578;
              heapClock = ~ heapClock;
        end

       2578 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1238] = 0;
              ip = 2579;
        end

       2579 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1238];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2580;
              heapClock = ~ heapClock;
        end

       2580 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2628;
        end

       2581 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2582;
        end

       2582 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[517];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 2;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2583;
              heapClock = ~ heapClock;
        end

       2583 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1239] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2584;
              heapClock = ~ heapClock;
        end

       2584 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[533] = localMem[1239] + 1;
              ip = 2585;
        end

       2585 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[524];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2586;
              heapClock = ~ heapClock;
        end

       2586 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1240] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2587;
              heapClock = ~ heapClock;
        end

       2587 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[534] = localMem[1240];
              ip = 2588;
        end

       2588 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[534];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = localMem[533];                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2589;
              heapClock = ~ heapClock;
        end

       2589 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1241] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2590;
              heapClock = ~ heapClock;
        end

       2590 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[535] = localMem[1241];
              ip = 2591;
        end

       2591 :
        begin                                                                   // jNe
          //$display("AAAA %4d %4d jNe", steps, ip);
              ip = localMem[535] != 0 ? 2599 : 2592;
        end

       2592 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2592");
        end

       2593 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2593");
        end

       2594 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2594");
        end

       2595 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2595");
        end

       2596 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
          // $display("Should not be executed  2596");
        end

       2597 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
          // $display("Should not be executed  2597");
        end

       2598 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
          // $display("Should not be executed  2598");
        end

       2599 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2600;
        end

       2600 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2601;
        end

       2601 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[536] = 0;
              ip = 2602;
        end

       2602 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2603;
        end

       2603 :
        begin                                                                   // jGe
          //$display("AAAA %4d %4d jGe", steps, ip);
              ip = localMem[536] >= 99 ? 2618 : 2604;
        end

       2604 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[535];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2605;
              heapClock = ~ heapClock;
        end

       2605 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1245] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2606;
              heapClock = ~ heapClock;
        end

       2606 :
        begin                                                                   // not
          //$display("AAAA %4d %4d not", steps, ip);
              localMem[537] = !localMem[1245];
              ip = 2607;
        end

       2607 :
        begin                                                                   // jTrue
          //$display("AAAA %4d %4d jTrue", steps, ip);
              ip = localMem[537] != 0 ? 2618 : 2608;
        end

       2608 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[535];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 6;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2609;
              heapClock = ~ heapClock;
        end

       2609 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1246] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2610;
              heapClock = ~ heapClock;
        end

       2610 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[538] = localMem[1246];
              ip = 2611;
        end

       2611 :
        begin                                                                   // movRead1
          //$display("AAAA %4d %4d movRead1", steps, ip);
              heapArray  = localMem[538];                                                  // Address of the item we wish to read from heap memory
              heapIndex  = 0;                                                  // Address of the item we wish to read from heap memory
              heapAction = `Read;                                           // Request a read, not a write
              ip = 2612;
              heapClock = ~ heapClock;
        end

       2612 :
        begin                                                                   // movRead2
          //$display("AAAA %4d %4d movRead2", steps, ip);
              localMem[1247] = heapOut;                                                     // Data retrieved from heap memory
              ip = 2613;
              heapClock = ~ heapClock;
        end

       2613 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[539] = localMem[1247];
              ip = 2614;
        end

       2614 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[535] = localMem[539];
              ip = 2615;
        end

       2615 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2616;
        end

       2616 :
        begin                                                                   // add
          //$display("AAAA %4d %4d add", steps, ip);
              localMem[536] = localMem[536] + 1;
              ip = 2617;
        end

       2617 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2602;
        end

       2618 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2619;
        end

       2619 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1248] = localMem[535];
              ip = 2620;
        end

       2620 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 0;                                                // Index of element to write to
              heapIn      = localMem[1248];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2621;
              heapClock = ~ heapClock;
        end

       2621 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1249] = 1;
              ip = 2622;
        end

       2622 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 1;                                                // Index of element to write to
              heapIn      = localMem[1249];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2623;
              heapClock = ~ heapClock;
        end

       2623 :
        begin                                                                   // mov
          //$display("AAAA %4d %4d mov", steps, ip);
              localMem[1250] = 0;
              ip = 2624;
        end

       2624 :
        begin                                                                   // movWrite1
          //$display("AAAA %4d %4d movWrite1", steps, ip);
              heapArray   = localMem[517];                                                // Array to write to
              heapIndex   = 2;                                                // Index of element to write to
              heapIn      = localMem[1250];                                                 // Data to write
              heapAction  = `Write;                                         // Request a write
              ip = 2625;
              heapClock = ~ heapClock;
        end

       2625 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2626;
        end

       2626 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2627;
        end

       2627 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2628;
        end

       2628 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2629;
        end

       2629 :
        begin                                                                   // jmp
          //$display("AAAA %4d %4d jmp", steps, ip);
              ip = 2505;
        end

       2630 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2630");
        end

       2631 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
          // $display("Should not be executed  2631");
        end

       2632 :
        begin                                                                   // label
          //$display("AAAA %4d %4d label", steps, ip);
              ip = 2633;
        end

       2633 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[517];
              ip = 2634;
              heapClock = ~ heapClock;
        end

       2634 :
        begin                                                                   // free
          //$display("AAAA %4d %4d free", steps, ip);
              heapAction = `Free;
              heapArray  = localMem[518];
              ip = 2635;
              heapClock = ~ heapClock;
        end

       2635 :
        begin                                                                   // tally
          //$display("AAAA %4d %4d tally", steps, ip);
            ip = 2636;
        end
      endcase
      success = outMem[0] == 1 && outMem[1] == 2 && outMem[2] == 3 && outMem[3] == 4 && outMem[4] == 5 && outMem[5] == 6 && outMem[6] == 7 && outMem[7] == 8 && outMem[8] == 9 && outMem[9] == 10 && outMem[10] == 11 && outMem[11] == 12 && outMem[12] == 13 && outMem[13] == 14 && outMem[14] == 15 && outMem[15] == 16 && outMem[16] == 17 && outMem[17] == 18 && outMem[18] == 19 && outMem[19] == 20 && outMem[20] == 21 && outMem[21] == 22 && outMem[22] == 23 && outMem[23] == 24 && outMem[24] == 25 && outMem[25] == 26 && outMem[26] == 27 && outMem[27] == 28 && outMem[28] == 29 && outMem[29] == 30 && outMem[30] == 31 && outMem[31] == 32 && outMem[32] == 33 && outMem[33] == 34 && outMem[34] == 35 && outMem[35] == 36 && outMem[36] == 37 && outMem[37] == 38 && outMem[38] == 39 && outMem[39] == 40 && outMem[40] == 41 && outMem[41] == 42 && outMem[42] == 43 && outMem[43] == 44 && outMem[44] == 45 && outMem[45] == 46 && outMem[46] == 47 && outMem[47] == 48 && outMem[48] == 49 && outMem[49] == 50 && outMem[50] == 51 && outMem[51] == 52 && outMem[52] == 53 && outMem[53] == 54 && outMem[54] == 55 && outMem[55] == 56 && outMem[56] == 57 && outMem[57] == 58 && outMem[58] == 59 && outMem[59] == 60 && outMem[60] == 61 && outMem[61] == 62 && outMem[62] == 63 && outMem[63] == 64 && outMem[64] == 65 && outMem[65] == 66 && outMem[66] == 67 && outMem[67] == 68 && outMem[68] == 69 && outMem[69] == 70 && outMem[70] == 71 && outMem[71] == 72 && outMem[72] == 73 && outMem[73] == 74 && outMem[74] == 75 && outMem[75] == 76 && outMem[76] == 77 && outMem[77] == 78 && outMem[78] == 79 && outMem[79] == 80 && outMem[80] == 81 && outMem[81] == 82 && outMem[82] == 83 && outMem[83] == 84 && outMem[84] == 85 && outMem[85] == 86 && outMem[86] == 87 && outMem[87] == 88 && outMem[88] == 89 && outMem[89] == 90 && outMem[90] == 91 && outMem[91] == 92 && outMem[92] == 93 && outMem[93] == 94 && outMem[94] == 95 && outMem[95] == 96 && outMem[96] == 97 && outMem[97] == 98 && outMem[98] == 99 && outMem[99] == 100 && outMem[100] == 101 && outMem[101] == 102 && outMem[102] == 103 && outMem[103] == 104 && outMem[104] == 105 && outMem[105] == 106 && outMem[106] == 107;
      steps = steps + 1;
      finished = steps >  67460;
    end
  end

endmodule
